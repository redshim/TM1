其他媒体|1591840687|zhidao_baidu|电脑/网络|ZHO|2015-01-02 12:22:01|"卡罗拉|k3|k4|买哪个车子比较合适|请教网友给指点"||http://zhidao.baidu.com/question/1303653602907494979.html?entry=qb_browse_default|2015-01-02
其他媒体|1613271864|wenwen_soso|生活家居|ZHO|2015-01-16 00:29:02|东风悦达起亚k3怎么视频放不出来|东风悦达起亚k3怎么视频放不出来 5|http://wenwen.soso.com/z/q622133911.htm?ch=wtk.title|2015-01-16
其他社区|1613828266|360wenda|已解决|ZHO|2015-01-16 11:03:02|我的卡装在联想乐檬 k3的手机上变2g...|不识别吧 你换个手机 或者换个卡卡 试试有些卡质量不好兼容不了送给回答者一份礼物送香吻 赠言：好帅的回答 楼主送上香吻一枚 以表诚挚谢意！ 00x用微信扫描二维码分享至好友和朋友圈分享到：检举 -->答答好搜问答团队最勤劳最可爱的答答5分钟前下面是答答童鞋给您的小建议 您看靠谱吗？初来乍到 弄错了您不要生气哦(*^__^*)答答小贴士|http://wenda.so.com/q/1421373414725107|2015-01-16
其他媒体|1613937315|hexun|滚动新闻 > 全部新闻|ZHO|2015-01-16 12:14:01|起亚K32015款现车出售 最高让利5000元【图】|　　海口行情近日 中国汽车消费网编辑从东风悦达起亚海南创亿4S店了解到 店内起亚K3现车出售 目前购车最高让利5000元。感兴趣的消费者可以进店了解详情 以下是2015款起亚K3的具体的报价表：海口地区起亚4s店最新价格：起亚K3报价表（2015-01-16）车型指导价销售价优惠情况现车情况起亚K3 2015款 1.6L MT GL10.28万9.78万0.5万有现车起亚K3 2015款 1.6L AT GL11.28万10.78万0.5万有现车起亚K3 2015款 1.6L AT GLS12.48万11.98万0.5万有现车起亚K3 2015款 1.6L AT DLX13.18万12.68万0.5万有现车起亚K3 2015款 1.6L AT Premium14.38万13.88万0.5万有现车起亚K3 2015款 1.8L AT Premium14.98万14.48万0.5万有现车中国汽车消费网制表　　起亚K3各地行情信息请关注：http://auto.315che.com/qiyak3/articles__43.htm　　更多同级别车型价格变动信息请关注：http://www.315che.com/hq/　　基本介绍：2015款K3的前中网颜色变更 后保险杠和排气管也经过了重新设计 DLX AT及以上车型配备了椭圆形的镀铬排气管。2015款K3还新增珍珠白这一可选车身颜色。中控面板位置的空调按钮增加镀铬装饰 车内引入了更多软性材料装饰。2015款K3的主要竞争对手还是目前市场上主流的紧凑型轿车 例如现代朗动、本田凌派、雪佛兰科鲁兹等。和竞争对手相比 丰富的配置和个性的造型是吸引不少消费者选择K3的因素。起亚K3 指导价： 10.28～14.98 万 品牌：起亚图片(共767 张)　　配置　　车吧　　报价　　口碑(共133 条)315che.com　　配置详解　　GL配备了主副驾驶座安全气囊、ABS+EBD、多功能方向盘上下调节、行车电脑显示屏、前座中央扶手、前雾灯、大灯高度可调、后视镜电动调节、后视镜加热、手动空调。　　GLS多了日间行车灯、后排杯架、后座中央扶手、座椅高低调节、真皮方向盘、电动天窗、无钥匙启动系统以及选装配置倒车视频影像、真皮座椅、腰部支撑调节、前排座椅电动调节、电动座椅记忆、座椅通风、GPS导航系统、蓝牙/车载电话等。　　DLX在GLS的基础上又多了EBD+EBA+ASR、真皮座椅、后座出风口和温度分区控制。　　Premium作为最高配 新增了后视镜电动折叠、后视镜记忆、氙气大灯、电动座椅记忆、前排座椅加热、座椅通风、前排座椅电动调节、腰部支撑调节、方向盘换挡、定速巡航、胎压监测装置。自动挡还可选装前/后排头部气囊(气帘)。　　注：中国汽车消费网 (www.315che.com) 提供的价格信息为编辑采集的及时信息 价格仅供参考 车市行情天天变 消费者如需购买相关车型 应该尽快与具体经销商电联或当面洽谈。另 文中引用图片和推荐经销商仅为资料信息 与价格信息来源无关。　　起亚K3榆林现车充足 购车最高优惠1.4万 榆林行情近日 中国汽车消费网编辑从东风悦达.起亚榆林经销商处了解到 现购东风悦达起亚k3可享1.4万现金优惠 目前店内现车销售。感兴趣的消费者可以进店了解详情 以下是2015款起亚K3的具体的报价表：榆林地区起亚4S店最新价格：起亚K3报价表（2015-01-13）车型指导价销售价优惠情况现车情况起亚K3 2015...查看　　2015款起亚K3优惠现金0.7万元 现车供应 广州行情近日 中国汽车消费网编辑从广州粤标汽车销售服务有限公司了解到 购买起亚K3可优惠7000元 店内有现车。感兴趣的消费者可以进店了解详情 以下是2015款起亚K3的具体的报价表：广州地区起亚4S店最新价格：起亚K3报价表（2015-01-13）车型指导价销售价优惠情况现车情况起亚K3 2015款 1.6L M...查看　　起亚K3优惠增至1万元 颜色可选现车充足 广州行情近日 中国汽车消费网编辑从广州地区东风悦达起亚经销商了解到 店内起亚K3现金优惠1万元 有现车在售。感兴趣的消费者可以进店了解详情 以下是2013款起亚K3的具体的报价表：广州地区起亚4S店最新价格：起亚K3报价表（2014-12-24）车型指导价销售价优惠情况现车情况起亚K3 2013款 1.6L MT ...查看　　起亚K3现金优惠1.2万 现车资源充足销售 南京行情近日 中国汽车消费网编辑获悉 南京金起汽车店内起亚K3现车销售 颜色可选 目前购车部分车型可优惠1.2万元 促销时间 2014.12.22-2014.12.26。感兴趣的消费者可以进店了解详情 以下是2013款起亚K3的具体的报价表：南京地区起亚4S店最新价格：起亚K3报价表（2014-12-22）车型指导...查看（责任编辑：HA002）|http://auto.hexun.com/2015-01-16/172449413.html|2015-01-16
其他媒体|1667163779|zhidao_baidu|电子数码|ZHO|2015-02-19 12:31:02|请教飞飞看电影听流行 丹拿bm6a mk1和mk3怎么选||http://zhidao.baidu.com/question/1447305648059709820.html?entry=qb_browse_default|2015-02-19
其他媒体|1696915137|tianya|音乐天地|ZHO|2015-03-11 01:11:02|[摇滚爵士]经典爵士歌曲（个人整理）|一、Jazzamor（爵士情人乐队）　　听的比较多的一个组合 基本每首曲子都不错 简单列出几个。这个组合的其他曲子也是很不错的 有首《tonight》百度是搜索不到的。可惜了。电脑里有jazzamor乐队的《lazy sunday afternoon》专辑 14首都不错 喜欢就跟我要吧。　　1、《fly me to the moon》：　　http://mag.china.com.cn/online/huayangshengnian/02/bg.mp3　　2、《Lovin’ You》：　　http://file.saycupid.com/filedata/filestore7/clubdata/********/Jazzamor%20[A%20Piece%20Of%20My%20Heart]%20-%2010%20Lovin’%20You.wma　　3、《Einfach Leben》　　http://www.xr-vision.com/bg_music/music/Thecolorofyou.wma　　4、《Beautiful day》　　http://www.magzone.com/upload/online/yue30/yue/music1.mp3　　二、小野丽莎 　　声线不错 某国首席 Bossa Nova 女王 有不少经典作品。她的《moon river》也是不错的 百度搜不到。　　1、《La Vie En Rose 》玫瑰人生 　　http://kogshgd.com/mail/meiguirensheng.wma　　一首法国老歌 小野丽莎的经典代表作。　　2、《cachito》 　　http://www.xfxt.com.cn/xiaonei/Cachito.wma 　　3、《she wore a yellow ribbon》　　http://www.minwt.com/kiki/mp3/YouAreMySunshine.mp3　　4、《my boy》　　http://www.sk360.cn/flash/11.mp3　　5、《pretty world》　　http://www.fish-photo.com/fish-photo/music/%C7%E9%D4%B5.mp3《pikake》5、　　6、《sabah wu masa》　　http://www.sh-thg.com/thg_ad/bgsound.mp3　　三、 Nat King Cole  纳京高 　　|http://bbs.tianya.cn/post-music-157048-1.shtml|2015-03-11
其他媒体|1701693133|zhidao_baidu|生活|ZHO|2015-03-13 19:31:01|东风悦达起亚k3后排座椅怎样拆除||http://zhidao.baidu.com/question/1797080351272132867.html?entry=qb_browse_default|2015-03-13
其他媒体|1706296899|zhidao_baidu|生活|ZHO|2015-03-17 01:27:36|起亚k3丰田卡罗拉雪佛兰新科鲁兹那款好一下||http://zhidao.baidu.com/question/1511635055094385140.html?entry=qb_browse_default|2015-03-17
其他媒体|1706803898|zhidao_baidu|电脑/网络|ZHO|2015-03-17 11:13:01|东风日产轩逸和k3哪个舒适度好点||http://zhidao.baidu.com/question/1703954997937674980.html?entry=qb_browse_default|2015-03-17
其他媒体|1706803927|zhidao_baidu|电脑/网络|ZHO|2015-03-17 11:13:01|东风日产轩逸和k3哪个舒适度好点||http://zhidao.baidu.com/question/682239186913206492.html?entry=qb_browse_default|2015-03-17
其他媒体|1710234891|webcars|降价信息|ZHO|2015-03-19 09:57:01|[郑州]  起亚K3S最高现金优惠2.00万元 现车充足|"　　【万车网 郑州行情】近日 万车网郑州站编辑从东风悦达起亚河南广发4S店了解到 购起亚K3S最高现金优惠2.00万元 现车充足 颜色可选 感兴趣的朋友可与经销商联系。具体优惠信息请见下表：　　近期火爆活动：　　【全城最低价 组团买新车】万车网团车活动火爆进行中（点击进入）　起亚K3S郑州地区行情车型指导价（万元）经销商报价（万元）优惠幅度（万元）2014款 1.6L 手动GL10.188.60↘1.582014款 1.6L 自动GL11.189.60↘1.582014款 1.6L 手动GLS11.489.90↘1.582014款 1.6L 自动GLS12.4810.90↘1.582014款 1.6L 自动DLX13.1811.60↘1.582014款 1.6L 自动Premium14.3812.38↘2.002015年3月19日行情 车辆价格随时变动 敬请关注当地市场http://www.webcars.com.cn/万车网制表您询问和购车时说明您是""万车网用户"" 会得到更好的服务！《点击可查看郑州地区起亚4S店》　　与K3不同 起亚K3S前进气格栅尺寸明显缩小 前保险杠采用大嘴式设计 整车设计更加年轻动感。车身尺寸方面 起亚K3S长宽高分别为4365/1780/1460mm 轴距达到2700mm。车身颜色方面 起亚K3S有透明白、钻石银、檀木黑、暗樱红、汉玉白、钛银色和新雅蓝共7款车身颜色可选。【起亚K3S 外观】【起亚K3S 外观】　　内饰方面 起亚K3S与K3整体内饰布局保持高度一致 中控台采用不对称式设计 在搭配黑色仿碳纤维装饰后 车内驾驶氛围凸显运动气息。内饰配色方面 起亚K3S还增加了黑棕配色方案供消费者选择。配置方面 起亚K3S全系标配后扰流板、随速感应自动落锁、带有CD(MP3)+AUX+USB+iPod读取功能的音响系统、前排座椅安全带高度可调、前排电子预紧式安全带等配置。除入门级车型外 余下5款车型均配有倒车雷达。【起亚K3S 内饰】【起亚K3S 内饰】　　动力方面 起亚K3S搭载了1.6L自然吸气发动机 该发动机的最大功率为128马力 峰值扭矩为156N·m。传动方面 与之匹配的是6速手动或6速自动变速箱。　　经销商信息：　　东风悦达起亚河南广发起亚专营店　　地址：郑州市西三环与化工路交叉口向北1000米 路西(西环汽车公园内)　　销售热线：0371—********　　声明：　　本文中涉及到的车型价格为万车网编辑在经销商处采集到的真实当日价格。由于汽车价格经常变化 并且为单一经销商的个体行为 所以价格仅供参考。具体价格请您致电或到店与经销商详细商谈。文中图片为车型实拍图 价格信息与图片拍摄地点无关。    本文导航         责任编辑：关鑫  关键词：起亚K3S 东风悦达起亚 郑州悦达起亚 起亚k3 福瑞迪 起亚k5 起亚k2 起亚智跑 起亚k3s 起亚狮跑东风悦达起亚 K3S K3 河南广发       查看车型   实时报价  参数配置  实拍图片  热点资讯  评分评论  万车知道"|http://www.webcars.com.cn/review/20150319/106313.html|2015-03-19
其他媒体|1710443371|pingxiaow|新闻滚动|ZHO|2015-03-19 12:12:02|电影飓风营救3好看吗？电影飓风营救3影评及剧情介绍|电影飓风营救3好看吗？电影飓风营救3影评及剧情介绍2015-03-19 11:08:50  来源：深窗综合  责任编辑：评校网  网友评论 当页面出现错位（表格引起的错位）或内容显示不完整时候 请点击这里阅读全文 导演: 奥利维尔·米加顿 编剧: 吕克·贝松 / 罗伯特·马克·卡门 主演: 连姆·尼森 / 福里斯特·惠特克 / 法米克·詹森 / 玛姬·格蕾斯 / 多格雷·斯科特 / 萨姆·斯普卢尔 / 唐·哈维 / 丹兰·布鲁诺 / 勒兰德·奥瑟 / 大卫·沃肖夫斯基 / 强·格瑞斯 / 约翰尼·韦斯顿 / 安德鲁·博尔巴 / 朱迪·比彻 / 安德鲁·霍华德 类型: 动作 / 惊悚 / 犯罪 制片国家/地区: 法国 语言: 英语 / 俄语 上映日期: 2015-03-20(中国大陆) / 2014-12-16(柏林首映) / 2015-01-21(法国) 片长: 109分钟 又名: 即刻救援3(台) / 救参96小时3(港) / Tak3n 电影飓风营救3剧情介绍 前中情局探员布莱恩（连姆·尼森 Liam Neeson 饰）这次要拯救的不是被绑架的家人 而是他自己。布莱恩发现前妻遭受到残忍地杀害 自己竟被诬陷为杀妻的凶手。悲愤又失落的他为了洗刷冤屈 必须使出浑身解数 找出真相并揪出杀人凶手 同时还得躲避中情局、联邦调查局和警方的多方追缉；除此之外 更重要的任务 就是保护他身边唯一所剩并是最重要的亲人——他的女儿（玛姬·格蕾斯 Maggie Grace 饰）…… 以下是豆瓣电影对电影飓风营救3影评介绍 林文清：真不知道编剧把警察弄成这个样子是为了侮辱他们还是侮辱自己还是侮辱观众。。。每次看到那个黑胖探长又是握棋子又是缠皮筋一副我最智慧的样子我就被蠢得要心脏病发作…… 过客：话说在这一集中 救女儿将不再是主线。鼓掌！本片主要讲特工老爸的昔日搭档在一次特殊任务中全部卦挡 大叔意识到可能又有一个狂人要找他复仇 于是 大叔开始介入追查真相。他必须在有限的时间里查清楚 摆平一切 以免祸及家人。可随着案情的发展 一个当年不可告人的秘密浮出了水面 zykmilan：片头做得好惊艳！比2好在有更多伯恩的味道而不是一味打打杀杀救女儿/老婆。结尾小反转虽然并不高明但很讨喜。看在年过六十的连姆大叔还在玩命打 以及系列中这命途多舛的家庭（女儿被绑、老婆被绑、老婆被杀…我要哭了）的份上也得给好评啊。。。 更深的白色：只算能看。没有拯救的紧迫感是硬伤 而且从来不考虑collateral damage是价值观扭曲。导演太爱航拍了吧 而且最后追飞机boss战什么的标准环节都设计乏力 敷衍了事。 二货云：廉颇老矣 尚能饭也～看见连姆尼森一把年纪了还跳楼 砸垃圾桶 我的老腰都看疼了 不是救女不是救妻 这只是一个退休老特工的拼老命的复仇之路。。。而且还找到半路 都找错了仇家 大部分的恶斗主要是因为大叔不和警察合作闹出的事故 高速公路飙车造成的连带伤害真是无比巨大。。。。 安蓝·怪伯爵：这次不说演员只说编剧这两位~鸡贼如吕导儿10部完事儿名誉什么的盆满钵满了 “欧罗巴”玩儿命拍人贩都预订到6了 虽然很多都算不上太好的片 但至少看着够娱乐不装逼这不就足够了！另一位编剧罗伯特几乎包办了贝松所有系列电影剧本 也是够拼的 勇气可嘉！下一集后爹出狱又要祸害你闺女了吧大叔好累！ 殇潮 Icarus：感觉有些审美疲劳了。。。而且结尾很仓促 但看样子还能拍个4.。。。。最关心的其实是师　　评校网 详情请访问：http://www.pingxiaow.com/gundong/2015/0319/279946.html|http://www.pingxiaow.com/gundong/2015/0319/279946.html|2015-03-19
其他社区|1711107022|360wenda|待解决问题|ZHO|2015-03-19 19:31:03|东风悦达起亚-起亚k3手自一体的首付是多少 首付后每个月要付多|东风悦达起亚-起亚k3手自一体的首付是多少 首付后每个月要付多匿名网友分类： 购房置业被浏览13次10分钟前检举|http://wenda.haosou.com/q/1426760401725480|2015-03-19
其他媒体|1711348930|yoka|搭配日记|ZHO|2015-03-19 22:22:04|带上可爱的大天猫咪 大胆搭配新风尚！|"带上可爱的大天猫咪 大胆搭配新风尚！     4 0   阅读 回复      跳转到指定楼层      加关注   anacoppla   工作：货币：荣誉：住址：关注：粉丝：  帖子：152 精华：20注册时间：2012-10-25      [发消息][看主贴][只看该作者] 发表于 2015-3-19 21:21 1#   带上可爱的大天猫咪 大胆搭配新风尚！ Jilme面膜华丽套装|京东火热上市！ 迪奥梦幻美肌修颜乳 追求素颜无瑕美肌 赫莲娜神秘艳后睫毛膏 开启全新倾世之美 HR赫莲娜绿宝瓶「轻乳霜」 开启年轻美肤之旅 阿玛尼「黑钥匙」三宝 开启护肤新篇章  yoka社区             乍暖还寒的季节 保暖的同时穿出美丽优雅知性的女人味 是所有女性永远的追求。安娜今天和大家分享自己的搭配小心得呦。look1：黑色调搭配 红色调提亮不需要花枝招展 沉稳内敛的颜色是主色调 所以安娜选择了这件黑色的长呢大衣 简单的剪裁、经典的版型经久不衰。翻领设计干练精明 无论你去什么场合见什么人 这样的经典大衣总不会出错。这款大衣最出彩的地方 就是下摆立体红色的花朵 让衣服更加精致 女人就要如娇艳的花朵一般。      初春时节这样一顶羊毛呢帽是搭配首选 不论你是中分还是刘海、长发还是短发 都可以很好的驾驭它。帽檐的宽度适中 两侧稍留发髻可以起到很好的修饰脸型的作用 微微的荷叶形波浪衬托出优雅复古的气质。因为大衣是经典版型 所以搭配这样荷叶边的帽子是点睛之笔 这是属于自己的别致的优雅小细节。  一双美丽的高跟鞋是女人必不可少的。尖头视觉上拉长脚部线条 性感十足。细高跟干练利落 简约的设计更加大气 充满韵味。红色与衣服上的花朵相呼应 美美哒。  上身的颜色不宜过多 包包也选择了红色的 金属链条背带时尚感十足。    look2：棕色相互呼应成为经典 印花刺绣复古十足这套衣服更加日常休闲化 灰色呢子也是永不过时的经典 百搭又时尚。腰带的设计凸出女性的线条。亮点在于后背的刺绣设计 树枝上一只活灵活现的鹦鹉 周围点缀上一朵朵小花 可爱动人 充满了春天的生机。与众不同的后背的刺绣设计让你成为人海中的那个亮点。  棕色的雪地靴非常舒适哦。与其他雪地靴的单一颜色不同 安娜选择了有刺绣花朵的雪地靴与大衣相呼应 是不是非常特别的美呢。仅仅如此还不够 与棕色帽子成为首尾呼应哦！  再来张安娜非常喜欢的背部刺绣特写 非常精致的做工。  帽子也选择了棕色 安娜喜欢简约大方 颜色不能太多而且要有呼应哦。包包是渐变的咖啡条纹 方形小包配上这套衣服妥妥的。  look3：灰姑娘的蓝裙子 还有少不了水晶鞋当然啦 春天快要到了 不能缺少一些靓丽的色彩。最近超级火的《灰姑娘》给我带来无限灵感。这件泡泡袖的天蓝色毛衣温暖又舒适 宽松的设计给人带来一丝初春的慵懒气息、十分妩媚动人。湖蓝色的不规则大摆裙深得我心 飘逸灵动、不对称设计别出心裁十分吸引人的眼球。  仙气十足的一套搭配 不管是出街还是聚会 都是时尚时尚最时尚哦。配上银色高跟鞋闪亮夺目 鞋面的一个弧度的设计非常好看别有韵味 biling biling 走到哪里都是女神。衣服的设计感比较强、层次较多 所以搭配银色贝壳状小包 小巧玲珑也能衬托出这套仙气的衣服。是时候告别旧爱 迎接新气象啦 你的衣柜里需要几件“新面孔”。2015天猫新风尚 大胆爱新衣。微博：@AnaCoppla公共微信号：anacoppla私人微信：anacoppla007"|http://bbs.yoka.com/thread-7237791-1-1.html|2015-03-19
其他媒体|1789673609|zhidao_baidu|生活|ZHO|2015-05-08 09:41:02|起亚k3的发动机是一汽丰田卡罗拉淘汰下来的吗||http://zhidao.baidu.com/question/1176089271171861259.html?entry=qb_browse_default|2015-05-08
其他媒体|1848780405|zhidao_baidu|电脑/网络 > 硬件 > 显示器|ZHO|2015-06-11 21:03:02|k31.6gls和雷凌1.6家用选那个好在哪里|k31.6gls和雷凌1.6家用选那个好在哪里5 分钟前匿名分类：硬件来自：手机知道硬件|http://zhidao.baidu.com/question/490018385785782812.html?entry=qb_browse_default|2015-06-11
기타|1853763599|xda|三星Galaxy S III I9308 RSS|ZHO|2015-06-15 00:30:02|2015年山东移动营业员转聘试题 %答-案【+****-****】咨询包过|"[咨询求助]2015年山东移动营业员转聘试题 %答-案【+****-****】咨询包过[复制链接]  会计科会计科当前在线UID*******阅读权限10好友0帖子9精华0积分2注册时间2015-6-14最后登录2015-6-14门户文章0 精华0帖子9积分2 汉堡19 个注册时间2015-6-14发消息 发表于 57 秒前 显示全部楼层 阅读模式 注册个账号还能参加论坛各种活动哦~您需要 登录 才可以下载或查看 没有帐号？立即注册  x2015年山东移动营业员转聘试题 %答-案【+****-****】咨询包过( P9 b"" O/ D8 P+ R+ t 2015年山东移动营业员转聘考前时间及试题资料+卡卡****-**** V40 T  ?) a3 K9 K  m3 m1 l5 f: j  f- J* G; e2 O9 p4 A| j2 T 2015年山东移动营业员转聘考试【真题】+2015年山东移动营业员转聘考前时间及试题资料+****-****.(通过率100%)壹手打造.100%保证选 择我们=选 择成 功原题操作[诚信第一| 效率第一|考试大纲、考试真题、考试科目、考试资料4 ~"" E% a1 c& ~% w2 d- l6 q| A3 D2 o( @  G8 v' o' U9 L3 E; ]| L. c: Z/ Q; j| I& M) K# q  ^【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】6 [) ^7 U( v& v  ]8 H( J7 ?( u2 y* t/ R6 g$ Z7 ~【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】* c. y' x& ]4 d* m. A& p/ ]6 l: D4 o6 p* {% M' d9 p9 q& t/ z; s| C5 D6 K8 V5 m| k0 z0 {: M: ^% ]服 8 q8 H9 I0 [( t& {* [( Y( a! y- u  j4 e$ t4 d"" P0 Y【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】| @5 D; w9 G4 e% Y; r# Z"" z* U2 g$ d; A5 G4 i* N; l& r/ s/ m+ R9 ]8 c服 # H4 [5 R% z# D6 Q: S2 u4 L3 b6 z7 I' z# j【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】6 m"" l"" B' A4 Z0 E. }6 Q( r) B$ Q6 N$ {1 Z# j8 r& ^6 A5 O+ ?+ L# q服 ' M. g(  9 g# Y9 U5 s"" D! p# M+ e8 T- a' ~/ v) _& Q: j"" Q; O4 [4 Q+ f' c0 H' b| F3 S1 [* @ 2015年山东移动营业员转聘考试卷答题+「****-****.」& M6 ~9 Y6 n$ Y8 V# t) Q3 d0 \. Y  A# ]* [0 {9 t- v* }+ L| L' {/ W% f9 O: R 2015年山东移动营业员转聘考前时间及试题资料+****-****.(通过率100%)壹手打造.100%保证选 择我们=选 择成 功原题操作[诚信第一| 效率第一|考试大纲、考试真题、考试科目、考试资料8 M& R. e% ^2 C. s) P- ?2 Y: \$ S*  3 ?- v  {7 N. a| m5 ]- g"" s. {/ E 2015年山东移动营业员转聘考前时间及试题资料+****-****.考前试题有个小和尚 每天早上负责清扫寺庙院子里的落叶。清晨起床扫落叶实在是一件苦差事 尤其在秋冬之际 每一次起风时 树叶总随风飞舞落下。+****-****. +****-****. +****-****. +****-****.8 d& C8 G$ M5 O) `0 `' i每天早上都需要花费许多时间才能清扫完树叶 这让小和尚头痛不已。他一直想要找个好办法让自己轻松些。后来有个和尚跟他说：“你在明天打扫之前先用力摇树 把落叶统统摇下来 后天就可以不用扫落叶了。”$ Z. ^# M8 y* B6 t6 w* Q0 E; E% C"" i9 R* L# s5 y) N3 Q/ ~* Y; \+ e% i) J3 k6 f1 r. p! Q7 m; t7 K8 U& X0 O& p) }* \' g: L* n$ `. r+ o7 f8 i4 d* i+ @. M  x0 A; Q/  . [5 V' F: Q8 v( W 6 z"" z- l- M* u# ]$ {     ^* c& c' K| e3 v/ ^# v' I9 v+ g7 j1 @7 }0 j$ I. S1 j0 L; w! t& l) h小和尚觉得这是个好办法 于是隔天他起了个大早 使劲地猛摇树干 这样他就可以把今天跟明天的落叶一次扫干净了。一整天小和尚都非常开心。+ Q3 Z2 U6 N; F+ @* S8 A! U7 R+ B1 f. O4 X$ M% a9 C| z/ `. c9 i| n* P' o+ s3 o8 U7 d; ^: R- g3 r. x1 J  l3 C5 `| U- a2 o0 G$ H4 K2 v  H; P$ U3 i! e6 A% Z; [+ ^2 F| ^5 k5 v3 U: f0 K0 V8 F$ C5 {: i9 H  E. M0 D 1 S. k7 v1 U: A' {第二天 小和尚到院子一看 不禁傻眼了 院子里如往日一样落叶满地。9 K/ I"" d: `2 Z9 `- C: H7 _* ]+ R) }. x0 d/ G8 \! ]$ q1 u. m* n; f# N9 ?4 z: @$ F7 }5 b4 V8 i$ k; A2 n! ^2 A5 k  W3 L5 \6 i& w& z: F0 r7 l7 U"" W4 u3 Y: n# q8 U& n这时老和尚走了过来 对小和尚说：“傻孩子 无论你今天怎么用力 明天的落叶还是会飘下来。”小和尚终于明白了 世上有很多事是无法提前的 惟有认真地活好当下 才是最真实的人生态度。青山遮不住 毕竟东流去。该发生的你怎么阻挡也阻挡不了 不会发生的你再努力也没有用。把当下的事情做好了 就无怨无悔。9 ~% D$ X6 I( P| J; A5 W! D3 O& X* y+ A"" g"" d: x"" X4 ]( F0 [( `* z' d% l( \# K9 q! L9 z; [$ k1 t# }# u2 [8 I/ ]. \& y' B* R' ]; E1 M: n' }8 Z7 S2 S/ {' B: M- d$ X( P生活原本没有痛苦- S9 j. e8 W& g: J| E% h. I! ^7 h+ G8 K' ?| O9 m- u1 Y+ ^! L8 u* o$ P$ F"" `: H+ x1 w! B' j7 Y6 f- R1 {: y* z' ~' g0 v2 b- S# n; A8 ?6 Y. e  ^* f6  ! E+ H7 ]/ l& I3 n: Q) ~  l3 {0 _| }- I8 Z生活原本没有烦恼 当欲望之火被点燃后 烦恼就来敲你的心门了。* V* h( W/ f$ i* i. `; w. D6 s5 f. s0 R- h7 m"" P5 R' L. G- C"" D* M6 X( s"" u; o) k8 ^9 B"" q!  : o( F7 N# f7 R1 q3 a1 U1 J. f- S6 H0 h$ j9 g; v2 D# H( o ) u* r+ K7 Q| u3 P  d/ C. z# h- T6 n; i0 B* H& g* A! X: I8 g7 R| C生活原本没有痛苦 当你开始计较得失 贪求更多时 痛苦便来缠身了。+ k| a% f9 ]2 E8 }( n2 M9 u$ E! A+ e"" O& R0 A9 m| K. c$ B- r. F8 e2 K"" m' i# n$ A3 z5 Z' d9 m& ^1 l9 g: W( c& j& W+ a& Q+ C1 O# }- d' k7 T: @# i! J* U' N/ V# O"" n9 a1  : O: ]% } : g1 b* q& O# _/ K6 D$ t/ a"" }- H2 i: {: P5 N: a% f0 E7 v; o1 ~3 ?; z8 D| [4 m! a| q从前 有个百万富翁 每天让他劳神费心的事情跟他拥有的财富一样多。所以 他每天都愁眉紧锁 难得有个笑脸。6 L# X4 l| t+ @/ e( S; d- C. n- ]| ^* m5 ~3 w5 J  ]+ W2 I"" h5 ?) Q( ~2 @  T0 V0 ?7 f"" p6 N6 n& H7 q' z( E. L) A | Y( D# A; D/ {9 x$ Z0 r) _' s/ c. b: o"" L3 u% u"" X. C! J# [9 A: B4 B) ?百万富翁的隔壁 住着磨豆腐的小俩口。曾有谚语说 人生三大苦 打铁撑船磨豆腐。但磨豆腐的这小俩口却乐在其中 一天到晚歌声笑声逗圆梦乐声不断地传到百万富翁的家里。- P. c/ z$ e: T$ r/ l9 p8 s) R| i/ L7 }( t; o8 m"" q* ?* X! y/ a) ]6 z. ?! d3 q6 p: R! z7 Y1 ]* R7 [3 }$ ~' Y"" f- e. f( L2 Z- T9 m4 n3 M# u' A3 I: I! n- s1 r. e- t4 x1 T2 }9 W  N% \* i! a$ }& M# d5 c2 \' U 5 L( D1 D4 b! q/ i0 b; l# s. j7 ]0 \百万富翁的夫人问老公：“我们有这么多钱 怎么还不如隔壁家磨豆腐的小俩口快乐呢？”/ k. m9 r& e6 h$ U0 C- r$ ?* B) l7 ?# y2 s; z& A) t9 y5 P2 A! T( N6 v| c8 t$ Z) b% p8 w9 P| U4 f5 i! V0 V8 }! x  ` 0 i: T4 ["" h% q9 o& \3 _/ Q- b9 q+ m3 Y* @( F* S2 V* w& a"" q#  / _. ~5 K| Q: b5 l! L! A* u# R* h百万富翁说：“这有什么 我让他们明天就笑不出来。”5 e5 r: D' Q| u$ R1 G* K"" x* v) i* r. Y5 H; o5 I  Y6 j6 R) A8 U# k& l) \7 q- w. ?# n4 w. B| U| n0 }2 y"" }/ o$ Q5 ^! z& j( S$ H  n$ z' y7 M. C| K9 g3 j2 O* P. D/ b7 R+ c$ u/ b5 X* U& D到了晚上 百万富翁隔着墙扔了一锭金元宝过去。第二天 磨豆腐的小俩口果然鸦雀无声。原来这小俩口正在合计呢！他们捡到了天下掉下来的”金元宝后 觉得自己发财了 磨豆腐这种又苦又累的活儿以后是不能再做了。可是 做生意吧 赔了怎么办；不做生意吧 总有坐吃山空的一天。丈夫心里还想 生意要是做大了 是该讨房小的呢还是该休了现在这个黄脸婆；妻子则在琢磨 早知道能发财 当初就不该嫁给这臭磨豆腐的。寻思呀琢磨呀 之前快乐得很的小俩口现在谁也没有心思说笑了 烦恼已经开始占据他们的心。更令小俩口痛苦的是 为什么天上不能多掉几个金元宝呢 这样就能想买什么就买什么了啊？# w* D4 _+ D7 X8 D| `8 S"" Z# `4 ~/ N3 G: a- J# {+ [+ [4 o+ w- S* l: Y% z. O5 G"" X  u7 q' j+ {; L2 y5 T6 o. }% d6 h"" h' t1 x7 w: q/ _  Z. K4 t"" F& y+ l  J生活原本没有烦恼 当欲望之火被点燃后 烦恼就来敲你的心门了。0 V"" X+ N! M3 g0 ^"" f. O5 b. B( v| W7 e; p( j( b* F  `# Y* z) t; X; R| z0 S9 d; o( @+ {! f! Q9 A* b9 w9 d2 x' T+ v 8 K' v: {: ^| H0 v4 v% c| {; f$ Q| i; G( [# Q"" N8 R4  7 ?6 ^6 f  b; x3 l3 J9 z2 g. k0 x5 k( k5 p4 e生活原本没有痛苦 当你开始计较得失 贪求更多时 痛苦便来缠身了。$ T5 h| N6 z9  3 z9 \$ _+ Y- h$ z( E"" \4 n6 ]/ e- @4 [6 q0 u+ c  r* l6 ]0 }9 M- c2 T2 }% R; P' {9 c8 ]$ e"" Y+ {: ?1 [* Q# w! P4 @1 F)  & }. J$ s: f; g& _( v9 ~) @0 H/ A' u4 Y7 [- ~6 D9 Y0 m8 A9 Z ! v  S* W% W. W* c! u"" R8 a# H( V/ _$ V% \+ O0 e5 W% `7  3 ^4 D青春很易逝 珍惜当下才能少些追悔“孩子 趁年轻 何不埋头苦干 以成就一番事业呢？”有位老人劝告一位少年。) Y; m: n7 @3 n$ l3 h; z6 a& t' g* H) p- C-  # h6 Q3 S  r% X2 E! {8 Z1 G3 d. z+ p5 a/ H3 u  ^  \. ^+ Y; C+ B8 X- D) J* F"" G) @; d2 ]1 W| T  o: v% g8 k. {7 v5 t* b7 v| P# w  W5 C: C6 V1 {  B( g8 Z8 ?1 m7 D$ {/ j: ~& Y( B: q4 n* n- v' _: ]1 J0 l"" p| O0 W' T$ }: O"" ]: {少年满不在乎地回答说：“何必那么急呢？我的青春年华才刚刚开始 时间有的是！再说 我的美好蓝图还未规划好呢！”“时间可不等人啊！”老人说 并把少年引到一个伸手不见五指的地下室里。“我什么也看不见啊！”少年说。! _% O- E: {( S; f# D8 t. {8 \' l' d% F; M5 I/ c4 ?8 \% u! W- z6 {0 ~- G: M- B- h- D1 q$ X1 X5 s. E; t5 u| o! h' P# B| D& h"" p5 I: u$ V$ F4 G9 V( N% _9 A; K$ @- H6 o' ^8 ?* W5 P! v# ]: m# H1 f* U: X) Q| x3 x4 k3 K3 r8 j) \+ ]/ }' `6 ]* q5 V老人擦亮一根火柴 对少年说：“趁火柴未熄 你在这地下室里随便选一件东西出去吧。”/ o/ H0 k- o; n& t/  . T"" P) i+ {| I+ K* e' O6 t0 @! i  n) h4 {( Y7 v9 _6 J0 q& w3 G9 Z9 h% z2 `1 ?| t3 y! V0 O. o1 C5 U( K$ {  P# W1 D& Y) O% f2  9 H+ [2 b"" e/ f * e' o6 _2 `1 `/ k+ x少年借助微弱的亮光 四处努力辨认地下室的物品 还未等他找到一样东西 火柴就燃尽了 地下室顿时又变得漆黑一团。“我什么也没拿到 火柴就灭了！”少年抱怨道。7 d9 @9 j"" d7 W$ m/ _3 H# l/ s: [* V9 {1 h: }1 X. i: {* S2 J"" M$ P; `; ?% Z3 h# i! b7 P( c7 C4 V"" o/ \"" l& u$ H% e5 E1 L; F1 X7 L7 S/ d"" O6 t! d4 a' u; E( \"" M' `3 ~* g- O. o4 T: l0 U8 q% C1 c| ~% c+ Y) p : ^) l8 f; X| Q  K% q# G"" y2 E2 S& {& l4 n8 j3 \3 \. \* v. j老人说：“你的青春年华就如同这燃烧的火柴 转瞬即逝 朋友 你要珍惜啊！”"" t"" Y* R- A3 R6 U/ D& f+ c. v0 Z% {% {2 R- H& a  x0 l! Y/ k& i| e! S+ G. i/ e9 ^0 S1 [+ d3 D1 }/ l3 C- l% x6 p+ ^+ }8 X2 C) x3 B   s- Y0 g"" m( H/ G! P! \5 t"" U0 A8 ?* X2 a) Z| J* L9  & C( R| {$ I& _( q. y4 ~$ d| H  k  Y| D人生说短不短 长寿者亦能活到百岁；说长不长 弹指一挥间。只是 青山遮不住 毕竟东流去 若是待走到生命的终点 才后悔所走过的人生 就为时已晚了。与其到那时后悔 不如今天多做一点 至少回首的时候苦乐参半 眼泪与笑脸并存。少一分遗憾 就多了一分回味。9 z4 Y| ]6 ~5 K|  4 q+ J& F2 T0 U: F7 I8 C  y* E- u8 h/ g+ f- Y  V& j2 M+ t# D# O6 A2 U8 O| h% h% i% q/ d$ m6 }5 ?| K5 i& ^"" n! e0 z1 J% ~6 L( }  h & I# q2 n7 R3 }# E* ~0 E2 a9 c% b- P) X1 o1 j2 _8 _2 G: n. h2 L9 x7 [:  * w0 N) q* Z* \1 k苦难很肥沃 滋润人成长8 D6 ]$ j; s+ i2 z0 t$ [0 J) @0 e% g' O. g9 v' m6 J- V! u+ z5 Z  Z"" _. d| i% O5 B$ K"" @8 t3 q2 d3 y"" \3 M4 J"" H; ?% }- o* j  W7 `! g) }: z/ g4 N; @4 v1 O5 w; [& F- W6 M| D: z: T) C8 l"" T1 w降临到你身上的苦难 常常是上天要把你的心志磨励得得更加坚强 成长得更加更加挺拔。苦难对于一个乐意和迫切成长的人来说 是非常有营养的补品！% s#  "" i& u# h7 k. u' \& o+ l& H/ e/ s0 ~5 w3 b* x: m8  ' U- n+ a: _: q| F3 o5 N| W5 U& s' }; F; X| s9  / U1 c+ V"" j3 T2 v- M5 z7 ~5 e7 H4 l"" a  B1  ' T ' C0 n  ~#  / X0 i% y2 r: t. `. F* L3 e0 [8 a5 Q5 {1 a2 \7 n寒冬腊月 一个名为“滴水”的和尚去天龙寺拜见仪山禅师。外面下着很大的雪 可是仪山禅师却不让他进门。那个和尚就在门外一直跪着 这一跪就是三天。仪山的弟子看他可怜 纷纷为他求情。可是仪山说：“我这里不是收容所 不收留那些没有住处的人！”弟子们没有办法 只好纷纷走开。& x0 f+ ]2 M  u% r' v/ ~1 S- W2 W- r# ~* @/  7 W8 j% u+ s4 v. Z"" E6 M' x$ i+ S+ V2 f9 v7 x9 j: V  K; @( B( w# V1 j; r: K; @) X: {  A6 g1 ]9 j6 q1 g1 r  r- P; {4 q' h$ m5 V2 p. i+ [) z0 W( Z1 i+ l% G  p$  3 G5 ~( T) z4 d/ o7 z+ }: u5 j& h  L  m"" k7 Z到了第四天的时候 那个和尚身上皴裂的地方开始流血 他一次次地倒下又重新起来 但他依然跪在那里 雷打不动。仪山下令弟子：“谁也不准开门 否则就将他逐出门外！”1 \& w  ^4 D0 }0 d4 N- {  W$ u+ t/ R3 [; B' H6 V; m! V% M4 S; a6 U9 P/ L: L2 T) E9 L$ z4 M"" E; R"" `; J! G3 Y+ F| \) s* S0 W( a* O  l| X/ [) Q: o6 t# j/ B2 Z . S) o- ^/ A3 {% r$ C3 g( ~* L6 F; L: e7  + A2 Z( Q/ h! E  n. }( z( f' Y# u:  七天后 那个和尚支撑不住 倒了下去。仪山出来试了一下他的鼻子 尚且有一丝呼吸 于是便下令将他扶了进去。滴水终于进了仪山门下参学。+ ^4 s9 X3 ^! o.  | u% w# q% `| D& a) [  o' C& @( T& W* k; n5 b' W$ J+ x6 P. X1 p- l: y4 b2 m* C  S) S8 C' N) \  y: L! Y0 g; X* U0 _. T: G& a2 q8 a* l8 w7 H% B. V; J| ]"" j1 B2 U; p' m| I/ Q4 D* M0 e"" p/ [+ E/  ( N * l1 g3 v/ L2 U; F$ y"" t$ Q3 j/ _有一天 滴水和尚向仪山禅师问道：“无字 与般若有什么分别？”& U% f2 ]: R; r4 q% w$ d0 @% \; d4 S/ [5 B- B  C: Z0 _0 }5 f; I. H3 k: }( O4 e. D( X! m3 H1 v; P/ H$ `3 N8 ^# q"" q# W4 o* [8 D. X- f9 l- r. o& z+ L. d6 G' R9 c2 K) }8 q"" X/ B1 B+ `: u' J* f/ U5 ]& R5 C2 Y8 ?6 `"" F! Y! J0 z$ P8 @话刚说完 仪山就一拳打了过来 并大吼道这个问题岂是你能问的？滚出去！”)  ' Q! T9 V. h: H$ W; a* U| s6 O7 W( s0 A. Y% K' b/ E% ^2 x"" x- L7 n+ {) V4 @2 R- N9 z8 q6 M- u; B' K# q7 h  d+ r$ H"" i! \( C/ ~( _ ' t  ^. P9 u+ c) Q"" O|  9 n7 Z) I: b% w) r9 M8  * f' j) K# U6 h滴水被仪山的拳头打得头晕目眩 耳朵里只有仪山的吼声 忽然间 滴水想通了：“有与无都是自己的肤浅意识 你看我有 我看我无。”  [$ s8 E8 A7 d3 w+ h! H! x: l0 _4 M) H5 ]   * g$ J"" s3 x! o# z1 j$ k| o: c2 T. U8 \- Z: P7 e# K- F6 }% h1 M2 ?) U 1 O1 a9 q* p& {' y- P. R0 q) N7 Y) C+ h5 v  z$ K. M4 ]- S* w0 i  j8 l"" ]5 ]  X$ ?( V# A0 K* U$ \9 b& F  C% T( ?- X还有一次 滴水感冒了 正在用纸擦鼻涕的时候 被仪山看到了 仪山大声喝道：“你的鼻子比别人的血汗珍贵？你这不是在糟蹋白纸吗？”滴水便不敢再擦了。4 ?* L) @5 @  w' l. J; Z6 p+ p$ U/ p& l5 x9 _( F( l  D5 q! g| ?| v9 W5 S; j6 [) c# C& J: x| A8 B8 s' ]6 w6 L! q/ q) W6 d. Q9 W* X2 C-  + i/ ^+ @# [2 ? 2 n0  & C+ i6 {. _& v1 P.  : K) c. T  m很多人都难以忍受仪山的冷峻 可滴水却说：“人间有三种出家人 下等僧利用师门的影响力 发扬光大自己；中等僧欣赏家师的慈悲 步步追随；上等僧在师父的键锤下日益强壮 终于找到自己的天空。”"" r2 T+ s! x# s6 L; O( e/ j# S& i* t; @3 J7 r! \6 H( e9 [0 T& f- O1  # x$ q& G: l$ W: T8 o7 p* x6 H( }'  ! y. z$ Z! @7 \/ C$ ^# O| V"" K/ A: A* t . W5 [& r7 c2 i5 R4 @- R* K) k( q7 m8 I+ N/  # x# Y9 M滴水和尚后来果然成为一代得道高僧。3 ]. x- `3 G"" o4 G| K% z7 h* q3 e8 t  [1 \: D+ Q( u|  0 B6 X( l| w4 s! E  w' v3 c; x. R8 p; K4 D: k"" }. \5 r/ B| R8 p/ Y# n| I5 K9 C2 `# v! K+ W     }5 D) o3 W8 z& G% D$ t( L( R/ z% D: U+ @9 ~+ T   1 G+ A1 r4 P! p1 s向你挥来的鞭子 常常是要你把头抬得更高 背脊挺得更直。4 [| x  F- Y"" z& u- x8 B* Y& N% a+ w| L2 p! m0 L9 }| z+ j5 B) C5 H6 p1 q/ w2 g  a& `) X* U+ X+ p"" O/ \3 z- n- q  E| w6 y9 N0 {: S# z% q7 M9 s5 \"" z! ?( j4 M9 ~| `3 p& q1 Z5 p+ m1 o1 V0 O6 \% k% q$ G' `/ j降临到你身上的苦难 常常是上天要把你的心志磨励得得更加坚强 成长得更加更加挺拔。苦难对于一个乐意和迫切成长的人来说 是非常有营养的补品！+ r* S+ N- J6 M' u9 W8 P' M$ N+ y! z- c/ l$ n) w5 w7 ?* X: o' x& A"" H/ @1 {1 r8 x; O3 U+ H  [2 E$  & V4 Q2 c/ ^# v: z  Q! b  W+ X( \' @ / _/ ^6 ^4 M) {| M8 b& K2 R. U# J3 H* W! @: x+ P) p* W' W; a/ b% I"" B6 S$ }& v7 L活出生命真意义. l( @* I5 ]& j  D9 Y) c0 u) g3 V% m' N3 w  H5 p0 F0 A: \; O; z* \* Z| I| I# A  d%  * @% b% v6 N- K7 ~6 U' E8 f0 S$ K"" r: q! N7 e* l# C* d* O- e4 }2 t6 Q; u9 Z% ]* b9 ?"" m5 w) e: q: M7 E 4 W0 V5 @"" w6 _; E( w% ~4 O: J$ D! j  n9 l1 Q2 `0  3 q) ~5 x6 E$ ?1 B# ?9 [6 e/ K$ ~' L/ M3 R: r$ Q% \7 n"" E| l4  . y& b' V. n; b4 j4 y0 R: ~! s"" c8 d* N+ B% f8 k( X : g) k  Y5 N$ S9 J6 w+ b& {$ \' B9 W0 Y& f( W5 A 8 T# n  }2 d2 K( R6 E| ~: U7 n( W& A) y3 D5 O3 [( t5 [6 {& z4 U& K! F% B; z; r/ h2 h| Z+ q# g0 o% H4 {4 c8 l3 l2 g/ q| F) {  Q* k1 `  a8 J1 c( Z4 L! g* r8 u* q; m$ E/ ~+ k: r / k! E/ t"" n1 \- g$ Z)  $ e7 @- W0 g7 \: o3 W5 k0 A1 a| r7 J( A; Y( n9 @0 L- ?"" j/ F# k+ i* N! J- s: V. [8 t. D0 P1 O( b2 Z ! j$ D. G- a! }( X4 m7 s2 ?! H& C& ~# Z) D: s1 u1 J% R! S7 k9 S | a/ O/ x+ D* w/ o9 v: b$ o   ! }. ~3 G: u5 a& l| R0 Z! v/ Q' L / T- e& X7 y1 t|  3 i; T. v8 M1  5 ~9 i  S 3 Z% G: E6 j"" v# ?"" V3 l: f5 U  z6 n5 N8 G| `| I7 x  B| y6 s% d. A5 J# o + n"" ~% Z& U! D7 [) B! W  d# `"" G3 c' h: M| L; r' V  f2 L) B 7 R9 {& J* n' j/ Z4 O; A8 ^% O; L& n"" e9 Q| ]| ~"" I0 D: J$ o0 x3 D3 l( E; V+ B | n: I6 G: c6 p; x: M) y; H  e. D' h6 E$ M6 M! g+ g8 P5 F|  "|http://bbs.xda.cn/thread-14997699-1-1.html|2015-06-15
其他媒体|1854792171|hexun|滚动新闻 > 全部新闻|ZHO|2015-06-15 16:20:02|起亚K3全能SUV配置参数最新资讯优惠 最新钜惠开售 低价狂降多少？|"　　悦达起亚作为起亚在华的合资品牌 K3成为东风悦达起亚旗下引入的第三款K系列车型 K3已经在成都车展亮相 其搭载了与现代朗动相同的动力系统 1.6L及1.8L发动机 并于2012年10月15日左右上市。　　声明：腾信店内现车充足颜色齐全！无须预定|当天来提车当天就可开这您的爱车回家！让您不一样的感觉 　　起亚K3车型最新价格变化报价车型　　厂商指导价　　(万元)　　优惠金额　　(万元)　　裸车价　　(万元)　　成交价　　(万元)　　赠送　　礼包现车情况起亚K3 2015款 1.6L 自动Premium14.38↓ 4询价10.*******需要预订起亚K3 2015款 1.6L 自动GLS12.48↓ 4询价8.*******　　现车充足　　(透明白)起亚K3 2015款 1.6L 自动GL11.28↓ 4询价7.*******　　现车充足　　(透明白)起亚K3 2015款 1.6L 自动DLX13.18↓ 4询价9.*******　　现车充足　　(透明白)起亚K3 2015款 1.6L 手动GLS11.48↓ 4询价7.*******　　现车充足　　(透明白、暗樱红)起亚K3 2015款 1.6L 手动GL10.28↓ 4询价6.*******　　现车充足　　(透明白)购车赠送豪华礼包：全车膜（进口）、地胶、脚垫、凉垫、把套、鸡皮、掸子、发动机护板、车身封釉、地盘封塑、后舱垫、行李架、脚踏板、前后保险杠、DVD导航、原厂导航、倒车影像、倒车雷达、真皮座椅、挡泥板2015年6月04日行情 车辆价格随时变动 敬请关注当地市场k3前脸24小时热线电话：*********** 李经理24小时热线电话：*********** 李经理k3尾灯24小时热线电话：*********** 李经理24小时热线电话：*********** 李经理　　声明：本公司于多家品牌4S店合作多年 现已因部分4S店未完成销售目标 特在此之际 所有车系均以低价冲量销售中 网上所报价格均为实际销售价格 无任何附加条件 请广大客户放心购买。　　北京腾信全体员工期待您的光临 您的满意是我们服务的宗旨！　　营业时间:周一至周日（8:30―17:30）　　《诚信企业》 《诚信营销》 《榜样企业》　　厂家直销 价格优惠 现车充足 颜色齐全 可走全国 全国联保！ 购车当天我们会为您提供正规发票 合格证 保养手册 信息表 使用说明书等齐全　　北京腾信汽车销售有限公司　　全面创新、求真务实　　以人为本、共创辉煌　　24小时销售电话：*********** 联系人；李经理以上信息仅供参考 具体优惠信息以到店核算为主。　　如系本站原创文章 转载请注明出处：汽车中国。（责任编辑：HN666）"|http://auto.hexun.com/2015-06-15/176739862.html|2015-06-15
기타|1854841843|xda|三星Galaxy S III I9308 RSS|ZHO|2015-06-15 16:49:01|2015年甘肃甘南藏族一万名试题100%及答-案【+****-****】咨询包过|"[咨询求助]2015年甘肃甘南藏族一万名试题100%及答-案【+****-****】咨询包过[复制链接]  特认同特认同当前离线UID*******阅读权限10好友0帖子27精华0积分5注册时间2015-6-15最后登录2015-6-15门户文章0 精华0帖子27积分5 汉堡56 个注册时间2015-6-15发消息 发表于 13 小时前 显示全部楼层 阅读模式 注册个账号还能参加论坛各种活动哦~您需要 登录 才可以下载或查看 没有帐号？立即注册  x2015年甘肃甘南藏族一万名试题100%及答-案【+****-****】咨询包过* H' [2 k0 Q; A- q! D9 k 2015年甘肃甘南藏族一万名考前时间及试题资料+卡卡****-**** V40 T  ?) a3 K9 K  m3 m1 l5 f: j  f9 c( [5 ^"" D( f;  5 @+ R 2015年甘肃甘南藏族一万名考试【真题】+2015年甘肃甘南藏族一万名考前时间及试题资料+****-****.(通过率100%)壹手打造.100%保证选 择我们=选 择成 功原题操作[诚信第一| 效率第一|考试大纲、考试真题、考试科目、考试资料4 ~"" E% a1 c& ~% w2 d- l6 q| A3 D2 o( @  G8 v' o' U9 L3 E; ]| L. c: Z% s: F2 f: b6 O% E1 w# M【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】6 [) ^7 U( v& v  ]8 H( J7 ?| W  I3 K; k"" A7 M: O; j【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】* c. y' x& ]4 d* m. A& p/ ]6 l: D4 o6 p* {% M' d9 p9 q& t/ z; s| C5 D# a4 _- p2 N: u服 8 q8 H9 I0 [( t& {* [( Y5 w6 [# ~/ H) H5 ?【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】| @5 D; w9 G4 e% Y; r# Z"" z* U2 g$ d; A5 G4 i* N: w' _# X7 T* o  m8 C; K服 # H4 [5 R% z# D6 Q: S% g0 y4 N5 d| ^5 d3 W1 u【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】 【+****-****.】6 m"" l"" B' A4 Z0 E. }6 Q( r) B$ Q6 N$ {1 Z# j| S/  | t% F$ l- C1 H服 ' M. g(  9 g# Y9 U5 s"" D! p# M+ e8 T- a' ~/ v) _& Q: j"" Q; O4 ["" o1 `| s6 M9 o& `0 v7 s 2015年甘肃甘南藏族一万名考试卷答题+「****-****.」& M6 ~9 Y6 n$ Y8 V# t) Q3 d0 \. Y  A# ]* [0 {9 t- v7 R"" C4 F) c9 Z0 `+ i5 o 2015年甘肃甘南藏族一万名考前时间及试题资料+****-****.(通过率100%)壹手打造.100%保证选 择我们=选 择成 功原题操作[诚信第一| 效率第一|考试大纲、考试真题、考试科目、考试资料8 M& R. e% ^2 C. s) P- ?2 Y: \$ S*  3 ?- v  {7 N. a| m0 {"" A3 H/ z( q6 M( y0 V| ?  D9 L 2015年甘肃甘南藏族一万名考前时间及试题资料+****-****.考前试题有个小和尚 每天早上负责清扫寺庙院子里的落叶。清晨起床扫落叶实在是一件苦差事 尤其在秋冬之际 每一次起风时 树叶总随风飞舞落下。+****-****. +****-****. +****-****. +****-****.! X$ a$ L: i2  ( L# g9 L' k每天早上都需要花费许多时间才能清扫完树叶 这让小和尚头痛不已。他一直想要找个好办法让自己轻松些。后来有个和尚跟他说：“你在明天打扫之前先用力摇树 把落叶统统摇下来 后天就可以不用扫落叶了。”$ Z. ^# M8 y* B6 t6 w* Q0 E; E% C"" i9 R* L# s5 y) N3 Q/ ~* Y; \+ e% i) J3 k6 f1 r. p! Q7 m; t7 K8 U& X0 O& p) }* \' g: L* n$ `. r+ o7 f8 i4 d* i+ @. M  x0 A; Q/  ' y; W4 ?5 j$ \- _- w5 ?' d) E' H 6 z"" z- l- M* u# ]$ {     ^* c& c' K| e3 v/ ^# v' I9 v+ g7 j1 @7 }0 j$ I. S1 j0 L; w! t& l) h小和尚觉得这是个好办法 于是隔天他起了个大早 使劲地猛摇树干 这样他就可以把今天跟明天的落叶一次扫干净了。一整天小和尚都非常开心。+ Q3 Z2 U6 N; F+ @* S8 A! U7 R+ B1 f. O4 X$ M% a9 C| z/ `. c9 i| n* P' o+ s3 o8 U7 d; ^: R- g3 r. x1 J  l3 C5 `| U- a2 o0 G$ H4 K2 v  H; P$ U3 i! e6 A% Z; [+ ^2 F| ^5 k5 v3 U: f0 K0 V- a' u( \. Y! f2 d4 k- C. S4 \2 T4 Z 1 S. k7 v1 U: A' {第二天 小和尚到院子一看 不禁傻眼了 院子里如往日一样落叶满地。9 K/ I"" d: `2 Z9 `- C: H7 _* ]+ R) }. x0 d/ G8 \! ]$ q1 u. m* n; f# N9 ?4 z: @$ F7 }5 b4 V8 i$ k; A2 n! ^- u+ ["" A3 c; T:  0 r& w& w& z: F0 r7 l7 U"" W4 u3 Y: n# q8 U& n这时老和尚走了过来 对小和尚说：“傻孩子 无论你今天怎么用力 明天的落叶还是会飘下来。”小和尚终于明白了 世上有很多事是无法提前的 惟有认真地活好当下 才是最真实的人生态度。青山遮不住 毕竟东流去。该发生的你怎么阻挡也阻挡不了 不会发生的你再努力也没有用。把当下的事情做好了 就无怨无悔。9 ~% D$ X6 I( P| J; A5 W! D3 O& X* y+ A"" g"" d: x"" X4 ]( F0 [( `* z' d% l( \# K9 q! L9 z; [$ k1 t# }  ?"" \; G; `5 d* ]8 ]' ]; E1 M: n' }8 Z7 S2 S/ {' B: M- d$ X( P生活原本没有痛苦- S9 j. e8 W& g: J| E% h. I! ^7 h+ G8 K' ?| O9 m- u1 Y+ ^! L8 u* o$ P$ F"" `: H+ x1 w! B' j7 Y6 f$ [0 X' G7 z; l( ^% D; h0 v2 b- S# n; A8 ?6 Y. e  ^* f6  ! E+ H7 ]/ l& I3 n: Q) ~  l3 {0 _| }- I8 Z生活原本没有烦恼 当欲望之火被点燃后 烦恼就来敲你的心门了。* V* h( W/ f$ i* i. `; w. D6 s5 f. s0 R- h7 m"" P5 R' L. G- C"" D* M6 X( s"" u; o) k8 ^9 B"" q!  : o( F7 N# f7 R1 q3 a1 U1 J. f- S6 H0 h& Q( `* s5 a0 V8 ^1 P( T6 L ) u* r+ K7 Q| u3 P  d/ C. z# h- T6 n; i0 B* H& g* A! X: I8 g7 R| C生活原本没有痛苦 当你开始计较得失 贪求更多时 痛苦便来缠身了。+ k| a% f9 ]2 E8 }( n2 M9 u$ E! A+ e"" O& R0 A9 m| K. c$ B- r. F8 e2 K"" m' i# n$ A3 z5 Z' d9 m& ^1 l9 g: W( c& j& W+ a& Q+ C1 O# }- d' k7 T: @# i! J* U' N/ V6 V  E% d5 {) m. v2 \ : g1 b* q& O# _/ K6 D$ t/ a"" }- H2 i: {: P5 N: a% f0 E7 v; o1 ~3 ?; z8 D| [4 m! a| q从前 有个百万富翁 每天让他劳神费心的事情跟他拥有的财富一样多。所以 他每天都愁眉紧锁 难得有个笑脸。6 L# X4 l| t+ @/ e( S; d- C. n- ]| ^* m5 ~3 w5 J  ]+ W2 I"" h5 ?) Q( ~2 @  T0 V0 ?7 f"" p6 N6 n* }% J) {! o* i& } | Y( D# A; D/ {9 x$ Z0 r) _' s/ c. b: o"" L3 u% u"" X. C! J# [9 A: B4 B) ?百万富翁的隔壁 住着磨豆腐的小俩口。曾有谚语说 人生三大苦 打铁撑船磨豆腐。但磨豆腐的这小俩口却乐在其中 一天到晚歌声笑声逗圆梦乐声不断地传到百万富翁的家里。- P. c/ z$ e: T$ r/ l9 p8 s) R| i/ L7 }( t; o8 m"" q* ?* X! y/ a) ]6 z. ?! d3 q6 p: R! z7 Y1 ]* R7 [3 }$ ~' Y"" f- e. f( L2 Z- T9 m4 n3 M# u' A3 I: I! n- s1 r. e- t4 x1 T2 }9 W  N5 o3 O; i! _- s+ N: R3 p 5 L( D1 D4 b! q/ i0 b; l# s. j7 ]0 \百万富翁的夫人问老公：“我们有这么多钱 怎么还不如隔壁家磨豆腐的小俩口快乐呢？”/ k. m9 r& e6 h$ U0 C- r$ ?* B) l7 ?# y2 s; z& A) t9 y5 P2 A! T( N6 v| c8 t$ Z) b% p+ L3 h0 {0 ]- n* m- _ 0 i: T4 ["" h% q9 o& \3 _/ Q- b9 q+ m3 Y* @( F* S2 V* w& a"" q#  / _. ~5 K| Q: b5 l! L! A* u# R* h百万富翁说：“这有什么 我让他们明天就笑不出来。”5 e5 r: D' Q| u$ R1 G* K"" x* v) i* r. Y5 H; o5 I  Y6 j6 R) A8 U# k& l) \7 q- w. ?# n4 w. B| U| n0 }2 y) `0 p% o0 l. M5 u( I& j( S$ H  n$ z' y7 M. C| K9 g3 j2 O* P. D/ b7 R+ c$ u/ b5 X* U& D到了晚上 百万富翁隔着墙扔了一锭金元宝过去。第二天 磨豆腐的小俩口果然鸦雀无声。原来这小俩口正在合计呢！他们捡到了天下掉下来的”金元宝后 觉得自己发财了 磨豆腐这种又苦又累的活儿以后是不能再做了。可是 做生意吧 赔了怎么办；不做生意吧 总有坐吃山空的一天。丈夫心里还想 生意要是做大了 是该讨房小的呢还是该休了现在这个黄脸婆；妻子则在琢磨 早知道能发财 当初就不该嫁给这臭磨豆腐的。寻思呀琢磨呀 之前快乐得很的小俩口现在谁也没有心思说笑了 烦恼已经开始占据他们的心。更令小俩口痛苦的是 为什么天上不能多掉几个金元宝呢 这样就能想买什么就买什么了啊？# w* D4 _+ D7 X8 D| `8 S"" Z# `4 ~/ N3 G7 E/ Y% W1 o9 P* T* a# K0 F' X: Y% z. O5 G"" X  u7 q' j+ {; L2 y5 T6 o. }% d6 h"" h' t1 x7 w: q/ _  Z. K4 t"" F& y+ l  J生活原本没有烦恼 当欲望之火被点燃后 烦恼就来敲你的心门了。0 V"" X+ N! M3 g0 ^"" f. O5 b. B( v| W7 e; p( j( b* F  `# Y* z) t; X; R| z0 S9 d; o( @+ {! f! Q9 A* b7 I! \. I% u9 @0 ^; U( k/ y 8 K' v: {: ^| H0 v4 v% c| {; f$ Q| i; G( [# Q"" N8 R4  7 ?6 ^6 f  b; x3 l3 J9 z2 g. k0 x5 k( k5 p4 e生活原本没有痛苦 当你开始计较得失 贪求更多时 痛苦便来缠身了。$ T5 h| N6 z9  3 z9 \$ _+ Y- h$ z( E"" \4 n6 ]/ e- @4 [6 q0 u+ c  r* l6 ]0 }9 M- c2 T2 }% R; P' {9 c8 ]$ e"" Y+ {: ?1 [* Q# w! P4 @1 F)  & }. J$ s: f; g& _( v9 ~) @0 H/ A' u4 Y7 [3 J+ z% W7 [1 `( o- b1 g7 ~% x6 o ! v  S* W% W. W* c! u"" R8 a# H( V/ _$ V% \+ O0 e5 W% `7  3 ^4 D青春很易逝 珍惜当下才能少些追悔“孩子 趁年轻 何不埋头苦干 以成就一番事业呢？”有位老人劝告一位少年。) Y; m: n7 @3 n$ l3 h; z6 a& t' g* H) p- C-  # h6 Q3 S  r% X2 E! {8 Z1 G3 d. z+ p5 a/ H3 u  ^  \. ^+ Y; C+ B8 X- D) J* F"" G) @; d2 ]1 W| T  o: v% g8 k. {7 v5 t* b7 v| P# w  W5 C: C6 V1 {  B( g8 Z8 ?1 m7 D$ {/ j: ~& Y( B: q4 n* n- v' _: ]1 J: W$ _8 V2 G6 o9 b少年满不在乎地回答说：“何必那么急呢？我的青春年华才刚刚开始 时间有的是！再说 我的美好蓝图还未规划好呢！”“时间可不等人啊！”老人说 并把少年引到一个伸手不见五指的地下室里。“我什么也看不见啊！”少年说。! _% O- E: {( S; f# D8 t. {8 \' l' d% F; M5 I/ c4 ?8 \% u! W- z6 {0 ~- G: M- B- h- D1 q$ X1 X5 s. E; t5 u| o! h' P# B| D& h"" p5 I: u$ V$ F4 G9 V( N% _9 A; K$ @- H6 o' ^8 ?* W5 P! v# ]: m# H1 f* U: X/ A| S6 p5 [+ P% i; s| y8 j) \+ ]/ }' `6 ]* q5 V老人擦亮一根火柴 对少年说：“趁火柴未熄 你在这地下室里随便选一件东西出去吧。”/ o/ H0 k- o; n& t/  . T"" P) i+ {| I+ K* e' O6 t0 @! i  n) h4 {( Y7 v9 _6 J0 q& w3 G9 Z9 h% z2 `1 ?| t3 y! V0 O. o1 C5 U( K$ {- z3 f- x(  6 f/ z; ?8 E * e' o6 _2 `1 `/ k+ x少年借助微弱的亮光 四处努力辨认地下室的物品 还未等他找到一样东西 火柴就燃尽了 地下室顿时又变得漆黑一团。“我什么也没拿到 火柴就灭了！”少年抱怨道。7 d9 @9 j"" d7 W$ m/ _3 H# l/ s: [* V9 {1 h: }1 X. i: {* S2 J"" M$ P; `; ?% Z3 h# i! b7 P( c7 C4 V"" o/ \"" l& u$ H% e5 E1 L; F1 X7 L7 S/ d"" O6 t! d4 a' u; E( \"" M' `3 ~* g- O. o5 R. F| ~8 ]0 i"" V"" S3 R& Z : ^) l8 f; X| Q  K% q# G"" y2 E2 S& {& l4 n8 j3 \3 \. \* v. j老人说：“你的青春年华就如同这燃烧的火柴 转瞬即逝 朋友 你要珍惜啊！”"" t"" Y* R- A3 R6 U/ D& f+ c. v0 Z% {% {2 R- H& a  x0 l! Y/ k& i| e! S+ G. i/ e9 ^0 S1 [+ d3 D1 }/ l3 C- l% x( `3 ]$ d+ ?2 e6 K0 L) @   s- Y0 g"" m( H/ G! P! \5 t"" U0 A8 ?* X2 a) Z| J* L9  & C( R| {$ I& _( q. y4 ~$ d| H  k  Y| D人生说短不短 长寿者亦能活到百岁；说长不长 弹指一挥间。只是 青山遮不住 毕竟东流去 若是待走到生命的终点 才后悔所走过的人生 就为时已晚了。与其到那时后悔 不如今天多做一点 至少回首的时候苦乐参半 眼泪与笑脸并存。少一分遗憾 就多了一分回味。9 z4 Y| ]6 ~5 K|  4 q+ J& F2 T0 U: F7 I8 C  y* E- u8 h/ g+ f- Y  V& j2 M+ t# D# O6 A2 U8 O| h% h% i% q/ d$ m6 }5 ?| K5 i& ^"" n& ?0 U7 d. B: ^8 A7 p & I# q2 n7 R3 }# E* ~0 E2 a9 c% b- P) X1 o1 j2 _8 _2 G: n. h2 L9 x7 [:  * w0 N) q* Z* \1 k苦难很肥沃 滋润人成长8 D6 ]$ j; s+ i2 z0 t$ [0 J) @0 e% g' O. g9 v' m6 J- V! u+ z5 Z  Z"" _. d| i% O5 B$ K"" @8 t3 q2 d3 y"" \3 M4 J1 k) [| r- k0 V| l' [) }: z/ g4 N; @4 v1 O5 w; [& F- W6 M| D: z: T) C8 l"" T1 w降临到你身上的苦难 常常是上天要把你的心志磨励得得更加坚强 成长得更加更加挺拔。苦难对于一个乐意和迫切成长的人来说 是非常有营养的补品！% s#  "" i& u# h7 k. u' \& o+ l& H/ e/ s0 ~5 w3 b* x: m8  ' U- n+ a: _: q| F3 o5 N| W5 U& s' }; F; X| s9  / U1 c+ V"" j3 T2 v- M5 z7 ~5 e# x) O  D/ u  R ' C0 n  ~#  / X0 i% y2 r: t. `. F* L3 e0 [8 a5 Q5 {1 a2 \7 n寒冬腊月 一个名为“滴水”的和尚去天龙寺拜见仪山禅师。外面下着很大的雪 可是仪山禅师却不让他进门。那个和尚就在门外一直跪着 这一跪就是三天。仪山的弟子看他可怜 纷纷为他求情。可是仪山说：“我这里不是收容所 不收留那些没有住处的人！”弟子们没有办法 只好纷纷走开。& x0 f+ ]2 M  u% r' v/ ~1 S- W2 W- r# ~* @/  7 W8 j% u+ s4 v. Z"" E6 M' x$ i+ S+ V2 f9 v7 x9 j: V  K; @( B( w# V1 j; r: K; @) X: {  A6 g1 ]9 j6 q1 g1 r1 H$ r& ?' N2 m"" v) z0 W( Z1 i+ l% G  p$  3 G5 ~( T) z4 d/ o7 z+ }: u5 j& h  L  m"" k7 Z到了第四天的时候 那个和尚身上皴裂的地方开始流血 他一次次地倒下又重新起来 但他依然跪在那里 雷打不动。仪山下令弟子：“谁也不准开门 否则就将他逐出门外！”1 \& w  ^4 D0 }0 d4 N- {  W$ u+ t/ R3 [; B' H6 V; m! V% M4 S; a6 U9 P/ L: L2 T) E9 L$ z4 M"" E; R"" `; J! G3 Y+ F| \) s* S0 W( a* O  l| X# D$ M6 g! c. a) @' T"" c; T . S) o- ^/ A3 {% r$ C3 g( ~* L6 F; L: e7  + A2 Z( Q/ h! E  n. }( z( f' Y# u:  七天后 那个和尚支撑不住 倒了下去。仪山出来试了一下他的鼻子 尚且有一丝呼吸 于是便下令将他扶了进去。滴水终于进了仪山门下参学。+ ^4 s9 X3 ^! o.  | u% w# q% `| D& a) [  o' C& @( T& W* k; n5 b' W$ J+ x6 P. X1 p- l: y4 b2 m* C  S) S8 C' N) \  y: L! Y0 g; X* U0 _. T: G& a2 q8 a* l8 w7 H% B. V; J| ]"" j1 B2 U; p' m| I/ Q$ W7 d9 }* o! h1 P * l1 g3 v/ L2 U; F$ y"" t$ Q3 j/ _有一天 滴水和尚向仪山禅师问道：“无字 与般若有什么分别？”& U% f2 ]: R; r4 q% w$ d0 @% \; d4 S/ [5 B- B  C: Z0 _0 }5 f; I. H3 k: }( O4 e. D( X! m3 H1 v; P/ H$ `3 N8 ^# q"" q# W4 o* [8 D. X- f9 l- r. o& z+ L. d6 G' R9 c2 K) }8 q"" X/ B1 B+ `3 k* S/ `; k3 g  \2 Y8 ?6 `"" F! Y! J0 z$ P8 @话刚说完 仪山就一拳打了过来 并大吼道这个问题岂是你能问的？滚出去！”)  ' Q! T9 V. h: H$ W; a* U| s6 O7 W( s0 A. Y% K' b/ E% ^2 x"" x- L7 n+ {) V4 @2 R- N9 z8 q6 M- u; B' K# q7 h9 l| k7 d3 E4 F9 g7 r6 m4 o6 U"" ] ' t  ^. P9 u+ c) Q"" O|  9 n7 Z) I: b% w) r9 M8  * f' j) K# U6 h滴水被仪山的拳头打得头晕目眩 耳朵里只有仪山的吼声 忽然间 滴水想通了：“有与无都是自己的肤浅意识 你看我有 我看我无。”  [$ s8 E8 A7 d3 w+ h! H! x: l0 _4 M) H5 ]   * g$ J"" s3 x! o# z1 j$ k| o: c2 T. U8 \- Z: P3 i' f+ C0 m* y8 U 1 O1 a9 q* p& {' y- P. R0 q) N7 Y) C+ h5 v  z$ K. M4 ]- S* w0 i  j8 l"" ]5 ]  X$ ?( V# A0 K* U$ \9 b& F  C% T( ?- X还有一次 滴水感冒了 正在用纸擦鼻涕的时候 被仪山看到了 仪山大声喝道：“你的鼻子比别人的血汗珍贵？你这不是在糟蹋白纸吗？”滴水便不敢再擦了。4 ?* L) @5 @  w' l. J; Z6 p+ p$ U/ p& l5 x9 _( F( l  D5 q! g| ?| v9 W5 S; j6 [) c# C& J: x| A8 B8 s' ]6 w6 L! q/ q) W6 d4 j! ?5 U2 y"" { 2 n0  & C+ i6 {. _& v1 P.  : K) c. T  m很多人都难以忍受仪山的冷峻 可滴水却说：“人间有三种出家人 下等僧利用师门的影响力 发扬光大自己；中等僧欣赏家师的慈悲 步步追随；上等僧在师父的键锤下日益强壮 终于找到自己的天空。”"" r2 T+ s! x# s6 L; O( e/ j# S& i* t; @3 J7 r! \6 H( e9 [0 T& f- O1  # x$ q& G: l$ W: T8 o7 p* x6 H( }'  ! y. z$ Z! @7 \/ C$ ^( }/ A& H| u% ^% h* z . W5 [& r7 c2 i5 R4 @- R* K) k( q7 m8 I+ N/  # x# Y9 M滴水和尚后来果然成为一代得道高僧。3 ]. x- `3 G"" o4 G| K% z7 h* q3 e8 t  [1 \: D+ Q( u|  0 B6 X( l| w4 s! E  w' v3 c; x. R8 p; K4 D: k"" }. \5 r/ B| R8 p/ Y# n| I5 K9 C2 `# v! K+ W     }% P| s: I0 y. h. f+ q& W$ t( L( R/ z% D: U+ @9 ~+ T   1 G+ A1 r4 P! p1 s向你挥来的鞭子 常常是要你把头抬得更高 背脊挺得更直。4 [| x  F- Y"" z& u- x8 B* Y& N% a+ w| L2 p! m0 L9 }| z+ j5 B) C5 H6 p1 q/ w2 g  a& `) X* U+ X+ p"" O/ \3 z- n- q  E| w6 y9 N0 {: S# z% q3 Z4 S4 _0 V/ I7 }!  ! x! R+ P  X| `3 p& q1 Z5 p+ m1 o1 V0 O6 \% k% q$ G' `/ j降临到你身上的苦难 常常是上天要把你的心志磨励得得更加坚强 成长得更加更加挺拔。苦难对于一个乐意和迫切成长的人来说 是非常有营养的补品！+ r* S+ N- J6 M' u9 W8 P' M$ N+ y! z- c/ l$ n) w5 w7 ?* X: o' x& A"" H/ @1 {1 r8 x; O3 U+ H  [2 E$  & V4 Q3 U( c- L* J3 m) K  E / _/ ^6 ^4 M) {| M8 b& K2 R. U# J3 H* W! @: x+ P) p* W' W; a/ b% I"" B6 S$ }& v7 L活出生命真意义. l( @* I5 ]& j  D9 Y) c0 u) g3 V% m' N3 w  H5 p0 F0 A: \; O; z* \* Z| I| I# A  d%  * @% b% v6 N| M  c% J"" ]' `# @. g"" r: q! N7 e* l# C* d* O- e4 }2 t6 Q; u9 Z% ]* b9 ?"" m5 w) e: q: M7 E 4 W0 V5 @"" w6 _; E( w% ~4 O: J$ D! j  n9 l1 Q2 `0  3 q) ~5 x6 E$ ?1 B# ?9 [6 e/ K$ ~' L/ M3 R: r$ Q% \7 n"" E| l4  . y& b' V. n; b4 j4 y0 R: ~7 p) Z2 w+ b. e : g) k  Y5 N$ S9 J6 w+ b& {$ \' B9 W0 Y& f( W5 A 8 T# n  }2 d2 K( R6 E| ~: U7 n( W& A) y3 D5 O3 [( t5 [6 {& z4 U& K! F% B; z; r/ h2 h| Z+ q# g0 o% H4 {4 c8 l3 l2 g/ q| F) {  Q* k1 `  a8 J1 c( Z4 L2 d2 F1 V& ^% F8 E"" A"" h( n# @ / k! E/ t"" n1 \- g$ Z)  $ e7 @- W0 g7 \: o3 W5 k0 A1 a| r7 J( A; Y( n9 @0 L- ?"" j/ F# k+ i* N8 G$ I. `# u2 ]- d ! j$ D. G- a! }( X4 m7 s2 ?! H& C& ~# Z) D: s1 u1 J% R! S7 k9 S | a/ O/ x+ D* w/ o9 v: b$ o   ! }. ~3 G: Z7 n$ `: N( g7 M7 Q| A  D) X# y / T- e& X7 y1 t|  3 i; T. v8 M1  5 ~9 i  S 3 Z% G: E6 j"" v# ?"" V3 l: f5 U  z6 n5 N8 G| `| I7 C"" o0 w* W& c1 ? + n"" ~% Z& U! D7 [) B! W  d# `"" G3 c' h: M| L; r' V  f2 L) B 7 R9 {& J* n' j/ Z4 O; A8 ^% O; L& n"" e9 Q| ]| ~"" I0 D: }* z. Q. ]2 i. [ | n: I6 G: c6 p; x: M) y; H  e. D' h6 E$ M6 M! g+ g8 P5 F|  "|http://bbs.xda.cn/thread-14997796-1-1.html|2015-06-15
其他媒体|1854877998|zhidao_baidu|生活|ZHO|2015-06-15 17:10:02|"东风悦达起亚k31|6lglsa丁"|来自：手机知道江苏|http://zhidao.baidu.com/question/497646183679433324.html?entry=qb_browse_default|2015-06-15
其他媒体|1855206630|zhidao_baidu|电脑/网络 > 硬件 > 显示器|ZHO|2015-06-15 20:29:01|"想买台车|起亚k3|丰田卡罗拉|奔腾b50|大众宝来|福特新福克斯|哪款车值"|"想买台车|起亚k3|丰田卡罗拉|奔腾b50|大众宝来|福特新福克斯|哪款车值9 分钟前匿名分类：CPU来自：手机知道CPU"|http://zhidao.baidu.com/question/746275311482007652.html?entry=qb_browse_default|2015-06-15
其他媒体|1879753623|tianya|我爱购物|ZHO|2015-06-30 00:17:01|电视最便宜互联网电视风口到来(转载)|　　“就电视行业来看 无论从眼前还是长远来说 只有真正从用户需求上激发的创新力及体验力比拼才是电视企业最需要做的。”近日 中国电子商会副秘书长陆刃波对当前互联网电视行业竞争发展做出上述分析。　　纵观整个行业 在竞争已经白热化的电视市场 想要做从用户需求出发的“最好的电视”并不容易 除了乐视、小米风头正劲外 传统彩电品牌纷纷通过结盟阿里、腾讯移植互联网基因 而早期进入互联网电视领域的联想也带着“独立17TV”再次卷土重来。　　互联网电视新锐品牌酷开便不得不提 自从今年独立以来 酷开站在了互联网电视大发展的风口上 推出了多款独具特色、极具影响力的产品 从目前情况来看 其市场销量稳步提升 用户口碑也不断攀升 在小米、乐视等互联网品牌占据主要舆论的市场中 占得一席之地。　　酷开销量稳步提升　　今年4月1日 酷开独立后推出了首款融合年轻人、儿童、老人三个模式的电视机酷开A43以及配置更为高级55英寸大屏A55。　　其中A43以强悍的配置和亲民的1999元价格给互联网电视领域注入了新的活力：第一台融合三类人群使用模式、第一台主打亲情牌的互联网电视。引述酷开董事长王志国的话来说 正是因为酷开对用户体验的重视 才造就了如A43这样的产品。　　而据王志国微博透露 酷开还将于7月举行一场发布会。短短几个月的时间酷开便推出多款新品 其产品的研发速度和能力可见一斑。　　值得一提的是 刚刚过去的618大战中 尽管小米与乐视之间的口水战吸睛十足 但酷开也不甘示弱 4K U55、K50J及K49等产品一举夺得天猫、京东及苏宁易购等众多平台的销量第一 与小米、乐视一同晋身互联网电视的第一阵营。　　互联网企业用人之道　　脱离了创维的“呵护” 面对前有小米、乐视等互联网跨界厂商 后有海信、TCL和长虹等传统电视厂商的夹击 酷开在未来能否走的更扎实、更优异也颇具挑战性。目前 酷开产品的年销量仍维持在百万台级别 与传统电视厂商动辄千万台的销量却有差距 但王志国带领的酷开团队却给了公司未来发展更美好的遐想空间。　　从618期间小米与乐视的唇枪舌战 以及海信、酷开等厂商的加入便不难看出 当前电视市场互联网化将成大势所趋 互联网电视市场迎来百家争鸣的元年 在如此行业趋势面前 酷开具有良好的发展基础。　　作为一家互联网公司 酷开团队拥有开放、平等的互联网企业作风 扁平化的管理让每个人都有足够的发展空间 权利下放 大家的想法能够很好地落实。正如王志国所言 酷开轻松、开放的团队氛围 曾让创维集团很多人心生“羡慕” 都想参与进来。　　全面布局产品线　　诚然 小米与乐视等互联网企业拥有更多用户 互联网营销方式也更为娴熟 但在产品线布局方面却不如酷开、海信等品牌 小米目前仅有三款产品销售 而乐视也迟迟在消费者热衷的55寸4K如此重要的产品段上缺阵 难以满足不同用户的多维度需求。　　反观酷开 其拥有高端配置的U系列、极致性价比的K系列以及颠覆创新性的A系列三大产品线 涵盖低中高各价位 并从40英寸到65英寸全线覆盖 能够全方位满足消费者需求。　　尽管酷开已完全独立 但创维作为坚实的后盾 却赋予了酷开先天的优异性 目前酷开的生产仍依托创维 保证了产品的优良工艺及供货等问题 同时 不同于小米乐视的售后外包 酷开共享创维的售后体系 全国共有4950家门店 拥有6000名售后工程师可随时提供最高质的服务。不可否认 作为品牌保障 创维的支持背景足够强大。　　2015年互联网电视市场可谓是充满挑战与机遇 单飞的酷开虽然和众多创业公司一样面临着众多难题 但酷开得益于实力殷实的创维技术支持 以及自身能把握用户的真正需求 并保证产品研发速度、能力和销量的稳步上升 这些努力都使这家快速发展的公司面对挑战时变的更为从容。　　家庭影院品牌哪个好　　http://sqbijia.com/html/7/5/ 　　电视十大品牌　　http://sqbijia.com/html/7/1/ 　　空调那个牌子好　　http://sqbijia.com/html/7/2/ 　　音响优缺点　　http://sqbijia.com/html/7/7/ 　　DVD型号　　http://sqbijia.com/html/7/6/ 　　冰箱有哪些品牌　　http://sqbijia.com/html/7/3/ 　　海尔Haier 电视哪款性价比最高　　http://sqbijia.com/html/7/1/22.html　　熊猫PANDA 电视最便宜　　http://sqbijia.com/html/7/1/14.html　　海尔Haier 电视买什么好　　http://sqbijia.com/html/7/1/22.html　　松下PANASONIC 电视怎么用　　http://sqbijia.com/html/7/1/9.html　　京东方BOE 电视最便宜　　http://sqbijia.com/html/7/1/17.html　　乐华ROWA 电视好吗　　http://sqbijia.com/html/7/1/15.html　　清华同方THTF 电视怎么用　　http://sqbijia.com/html/7/1/12.html　　康佳KONKA 电视对比　　http://sqbijia.com/html/7/1/7.html　　夏普SHARP 电视选购　　http://sqbijia.com/html/7/1/1.html　　先锋 电视怎么用　　http://sqbijia.com/html/7/1/21.html　　东芝TOSHIBA 电视买什么好　　http://sqbijia.com/html/7/1/13.html　　TCL王牌 电视怎么样　　http://sqbijia.com/html/7/1/8.html　　http://www.haha2.com/tianya/p/768_511235.html　　http://wangxuzhi.diandian.com/post/2015-06-15/***********　　http://www.shuixiangu.com/thread-93882-1-1.html　　http://www.kx001.com/diary/view_*********_********.html　　http://********.blog.hexun.com/*********_d.html　　http://www.vapee.com/team/127645.html　　http://i.changturen.com/blog-10775-328.html　　http://www.tmallze.com/html/768_511235.html　　http://www.kx001.com/diary/view_*********_********.html　　http://www.0554.us/tianya/du/768_501727.html　　http://www.mywlyx.cn/thread-360934-1-1.html　　http://club.suohoo.com/thread-496060-1-1.html　　http://huaban.com/pins/*********/　　http://www.0554.us/tianya/du/768_509133.html　　http://bbs.ybtop.com/thread-792033-1-1.html　　http://t.qq.com/p/t/***************　　http://www.0554.us/tianya/du/768_499909.html　　http://www.shuixiangu.com/thread-93056-1-1.html　　http://www.0554.us/tianya/du/768_495025.html　　http://taoker.pintuxiu.com/detail-index-share_id-2671.html　　http://www.wealink.com/dangan/*******/　　http://liuningyuan.bokee.com/*********.html　　http://blog.cnfol.com/wanghxhx/article/1434******-*******89.html　　http://www.0554.us/tianya/du/768_502650.html　　http://blog.cnfol.com/wanghxhx/article/1435******-*******05.html　　http://www.0554.us/tianya/du/768_510000.html　　http://bbs.one120.com/2015-6/27/***********.html　　http://www.mywlyx.cn/thread-360439-1-1.html　　http://www.bbyz.com/blog/show_*******_198187.html　　http://blog.cnfol.com/wanghxhx/article/1434******-*******49.html　　http://blog.cnfol.com/wanghxhx/article/1434******-*******55.html　　http://www.tmallze.com/html/768_509133.html　　http://wangxuzhi.diandian.com/post/2015-06-25/***********　　http://wangxuzhi.diandian.com/post/2015-06-21/***********　　http://www.kktie.com/tieku/768_509992.html　　http://www.kktie.com/tieku/768_495025.html　　http://www.seee.com.cn/bbs/showtopic-********.aspx　　http://www.mywlyx.cn/thread-360138-1-1.html　　http://huaban.com/pins/*********/　　http://www.kktie.com/tieku/768_505732.html　　http://www.tmallze.com/html/768_505732.html　　http://www.shuixiangu.com/thread-93935-1-1.html　　http://www.shuixiangu.com/thread-92933-1-1.html　　http://www.ahmu.net/read.php?tid-150454-ds-1.html　　http://blog.cnfol.com/wanghxhx/article/1434******-*******31.html　　http://blog.cnfol.com/wanghxhx/article/1435******-*******77.html　　http://bbs.cz001.com.cn/read-htm-tid-*******.html　　http://blog.tianya.cn/post-5******-*******7-1.shtml　　http://www.tmallze.com/html/768_495025.html　　http://t.qq.com/p/t/***************　　http://blog.tianya.cn/post-5******-*******4-1.shtml　　http://********.blog.hexun.com/*********_d.html　　http://i.changturen.com/blog-10775-329.html　　http://bbs.cz001.com.cn/read-htm-tid-*******.html　　http://ziyouzizaiziyouziz.lofter.com/post/1d3e7065_7434d63/　　http://www.kktie.com/tieku/768_510000.html　　http://www.haha2.com/tianya/p/768_499909.html　　http://bbs.23qw.com/thread-294925-1-1.html　　http://www.vapee.com/team/127403.html　　http://weibo.com/p/******************2560　　http://www.vapee.com/team/127594.html　　http://www.shuixiangu.com/thread-93166-1-1.html　　http://bbs.ybtop.com/thread-793052-1-1.html　　http://www.tmallze.com/html/768_509992.html　　http://wenwen.sogou.com/z/q*********.htm　　http://blog.tianya.cn/post-5******-*******2-1.shtml　　http://www.kktie.com/tieku/768_503350.html　　http://show.sodao.com/show/*******　　http://weibo.com/p/******************9866　　http://bbs.23qw.com/thread-294927-1-1.html　　http://taoker.pintuxiu.com/detail-index-share_id-2667.html　　http://www.health720.com/info-id-*******.html　　http://bbs.one120.com/2015-6/28/***********.html　　http://tieba.baidu.com/p/**********　　http://www.health720.com/info-id-*******.html　　http://********.blog.hexun.com/*********_d.html　　http://t.qq.com/p/t/***************　　http://www.shuixiangu.com/thread-92776-1-1.html　　http://www.health720.com/info-id-*******.html　　http://********.blog.hexun.com/*********_d.html　　http://bbs.cz001.com.cn/read-htm-tid-*******.html　　http://www.vapee.com/team/127293.html　　http://www.tmallze.com/html/768_502650.html　　http://www.kktie.com/tieku/768_509133.html　　http://wenwen.sogou.com/z/q*********.htm　　http://www.bbyz.com/blog/show_*******_198186.html　　http://********.blog.hexun.com/*********_d.html　　http://www.tmallze.com/html/768_510000.html　　http://www.seee.com.cn/bbs/showtopic-********.aspx　　http://bbs.cz001.com.cn/read-htm-tid-*******.html　　http://liuningyuan.bokee.com/*********.html　　http://www.0554.us/tianya/du/768_505732.html　　http://taoker.pintuxiu.com/detail-index-share_id-2666.html　　http://www.docin.com/p-**********.html　　http://www.0554.us/tianya/du/768_503350.html　　http://weibo.com/p/********dcb73e60102vk3e　　http://wangxuzhi.diandian.com/post/2015-06-16/***********　　http://www.kktie.com/tieku/768_502650.html　　http://www.kktie.com/tieku/768_511235.html　　http://www.duitang.com/people/mblog/*********/detail/　　http://www.kktie.com/tieku/768_509118.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/5/484.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/5/255.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/6/2/9.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/2/25.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/11/51.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/10/1/19.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/7/7/31.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/7/8/4.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/3/290.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/5/270.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/2/314.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/4/28.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/6/1/59.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/13/29.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/1/2/82.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/1/2/48.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/2/9/7.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/11/6/15.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/1/2/46.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/10/13/17.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/3/9/22.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/9/115.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/2/199.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/10/10/41.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/11/21.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/4/6.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/7/10/24.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/3/1/48.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/11/187.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/6/41.html　　http://badlink.links.cn/?url=http://sqbijia.com/html/12/3/303.html|http://bbs.tianya.cn/post-768-512428-1.shtml|2015-06-30
其他社区|1881263545|360wenda|已解决|ZHO|2015-06-30 19:51:01|起亚k3有时路上打晃 是怎么回事？|"建议你检查下摆臂送给回答者一份礼物送香吻 赠言：好帅的回答 楼主送上香吻一枚 以表诚挚谢意！ 10x用微信扫描二维码分享至好友和朋友圈分享到：检举 -->答答好搜问答团队最勤劳最可爱的答答13分钟前下面是答答童鞋给您的小建议 您看靠谱吗？初来乍到 弄错了您不要生气哦(*^__^*)答答小贴士相关问题起亚K3后装的氙气大灯有时亮有时不亮的是怎么回事?22013.06.15起亚k3夏天开空调的时候油门踏板会变沉是怎么回事?不是发动...22014.07.10起亚K3日行灯开时|车后的小灯也要亮啊?是怎么回事?_12013.11.17起亚K2行驶一小段路发动机难冷却时怎么回事22014.10.06东风悦达起亚赛拉图车喇叭有时单音甚至无音|是怎么回事?2014.05.09查看更多关于的问题 >>"|http://wenda.haosou.com/q/1435660616616466|2015-06-30
其他媒体|1949726904|wenwen_sogou|生活家居|ZHO|2015-08-09 16:02:01|2013版东风悦达起亚k3手动高配带天窗车价能卖...|2013版东风悦达起亚k3手动高配带天窗车价能卖多钱？      补充：2013年8月买的|http://wenwen.sogou.com/z/q632349882.htm?ch=wtk.title|2015-08-09
其他媒体|1949899165|zhidao_baidu|生活|ZHO|2015-08-09 18:27:08|雷凌1.6手动低配跟k31.6手动低配哪个更适合购买|来自：手机知道汽车|http://zhidao.baidu.com/question/1605654298965516227.html?entry=qb_browse_default|2015-08-09
其他媒体|1973288881|zhidao_baidu|电子数码 > MP4/MP3|ZHO|2015-08-23 01:27:13|东风悦达起亚k3北京2手车多少钱|北京|http://zhidao.baidu.com/question/520943597473306325.html?fr=qlquick&entry=qb_list_default|2015-08-23
其他媒体|1973593057|zhidao_baidu|电脑/网络 > 电脑装机|ZHO|2015-08-23 09:49:01|东风悦达起亚k3左前车门下刮个窟窿可以修复吗|来自：手机知道汽车|http://zhidao.baidu.com/question/1496391129395559059.html?fr=qlquick&entry=qb_list_default|2015-08-23
其他媒体|1973846017|zhidao_baidu|电子数码 > 手机/通讯-手机使用|ZHO|2015-08-23 13:50:01|12年东风悦达起亚 k3 1.6 l 自动波箱油放油罗丝在什么位置|汽车|http://zhidao.baidu.com/question/362689205234286292.html?fr=qlquick&entry=qb_list_default|2015-08-23
其他媒体|1973895512|zhidao_baidu|生活 > 家电|ZHO|2015-08-23 14:36:01|马自达axela和k3和卡罗拉哪个好|汽车|http://zhidao.baidu.com/question/1692555751817616948.html?fr=qlquick&entry=qb_list_default|2015-08-23
其他媒体|1974568183|zhidao_baidu|游戏|ZHO|2015-08-23 23:29:01|东风悦达起亚k3得变速箱电脑版在那个位置?|来自：手机知道汽车东风悦达起亚k3得变速箱电脑版在那个位置?|http://zhidao.baidu.com/question/1576725680148940980.html?fr=qlquick&entry=qb_list_default|2015-08-23
其他媒体|2037213848|mobile01|新進文章|ZHO|2015-09-30 01:47:23|「Ford 好友默契出遊去」 kuga 2.0 柴油 台中到苗栗苑裡來回 優缺點|「Ford 好友默契出遊去」 fiesta 1.0 5D 台中到武嶺來回 優缺點台中高鐵站艾維士租車領車出發→74快速道路→國3高速公路→苗栗苑裡看熊貓彩繪稻田→國3高速公路→台中大雪山→台中艾維士還車路線包含平地、市區、爬坡、快速道路、高速公路、大雪山的山路等等最大馬力(ps/ rpm)	180 hp/3500 rpm最大扭力(kg-m/ rpm)	40.8 kgm/2000~2500 rpm車道偏移警示（LAS）、自動緊急煞車（SCBS）、主動巡航控制系統後座出風口+後座也可多衝手機充電也有藍色氣氛燈柴油版後座 有點+厚比汽油版好座一點點 比同級休旅車中 cx5 rav4 xtrail u6難坐了點 調整後座傾斜角度小了點 也有中間頭枕+中間後幅走 柴油版跟2.0汽油頂級旗艦版唯一10向電動可調座椅柴油版新引擎 180p 也比柴油所有休旅車更省油  舊款 focus mk3 163p mk3.5新馬丁頭 柴油 也改成180p 固特意牌 235-50-r18吋跑山路超穩定車道偏移警示超大天窗 只能開一半 不能開全部後車廂有平整化套件 伸縮後帳版沒備胎 有自動補胎劑後倒車攝影機 也會跟著自動轉彎出現綠色圖案 就是停紅燈會自動熄火 蛋也把冷氣給關閉 變成吹送風空調不想要自動熄火 左邊可按鈕 取消關閉 蛋每次發動 要自己多按鈕 高速公路 車道偏移 方向盤會震動 冷氣出風口沒銀色電鍍裝飾條不會有反光問題人跟好車-kuga 合照kuga優點表現好的地方1.隔音好 高速時有效隔絕風切聲 4門有上很多隔音條2.2.0柴油動力夠用 爬山路的波時油門輕踩輕鬆 在高速公路上開到160 底盤也很穩定3.跑山路測試懸吊表現Q彈比較舒適點 歐係車感覺4.全車系搭載ESP、ABS、EBD、EBA、斜坡起步輔助系統 除了 1.5 入門陽春2種款式 配5srs 全車系1.5+2.0汽油+2.0柴油標配7srs5.8顆喇叭sync系統 放mp3音樂音質也不錯 還有低音 中音 高音 可調7.左右後照鏡有廣角鏡片8.方向燈桿小壓一下閃3下9.駕駛座4個窗戶鍵 小案 全升上全升下10.開啟引擎蓋 裡頭有黃色超厚的保護殼 以免燙到手 11.爬陡坡放開煞車踏板會自動幫您煞住3秒免擔心會向後滑行！12.白天或晚上開車門也有照明燈亮起 開啟後車廂也會亮照明燈 按遙控器開啟厚車廂 前後左右方向燈會閃一下13.下雨天自動開啟雨刷快慢 雨刷配軟骨雨刷 開車不會被雨刷擋道視線14.進墜道自動開啟大燈！ 開啟大燈是圓形旋轉式跟日系車不一樣15.倒車時 有出現逼逼聲音 感應到旁邊有障礙物 音響播放音樂會自動關閉 專心避開障礙物 以免刮傷車子16.音響還在播放歌 引擎熄火後 開啟駕駛座車門 音響自動關閉17.關門聲很進口車關門感覺 不繪像日系車關上後都㕩 很大聲18.駕駛座挺類似賽車椅 有包覆性感覺19.18吋固特意牌輪胎跑高速公路上+山路還不錯21.右後座地板下方有小抽屜 可放女生用品缺點還需改善的地方1. 全車系沒配有視覺盲點偵測系統2.後座座椅椅背稍直 後座空間小了點 後座不夠厚也不夠長 傾斜角度不夠往後躺3.後座置物空間少 雜物無處放4.停紅燈自動熄火 採煞車 有時有出先自動熄火 有時沒自動熄火5.手動換檔系統建議還是更改到方向盤後撥片比較順6.自動熄火 自動關閉冷氣 改吹送風空調7.排n黨容易排到r黨8.大燈沒有魚眼+hid+led晝行燈 9.牌照燈沒有像focus 有白光的led 小燈也改led 也多增加led晝行燈 10.免費體驗開福特新車活動時沒有附上操作sync系統的說明書 需要摸索老半天才知道如何使用11.運動版能夠學focus 大燈有薰黑樣式12.按遙控開啟或關閉 只能從駕駛門打開 其他3個門鎖 沒開13.天窗很大 無法開啟全部 只能開一半14.厚照鏡摺疊收起 無法像focus和fiesta平整收全部 只能收一半15.沒胎壓偵測福特歐洲車 kuga 2.0 柴油渦輪版5D果然是台好車！感謝福特提供好友默契免費開新車出遊去充實的一天~|http://www.mobile01.com/topicdetail.php?f=260&t=4553909|2015-09-30
기타|2038548743|ngzb|新闻互动|ZHO|2015-09-30 19:28:02|建行开展信用卡境外消费促销活动 33万人次享受优惠|"马上注册 结交更多好友 享用更多功能 让你轻松玩转南宁您需要 登录 才可以下载或查看 没有帐号？立即注册  x建行龙卡信用卡遇“建”世界遇见你+ B"" _| v- [-  0 \! E) `* Z+ X　　今年上半年|我国出境旅游人次近6200万|每25人次中就有1人使用建设银行龙卡信用卡。建设银行开展信用卡境外消费促销活动一年来|已有33万人次的客户享受了境外线上及线下优惠。想成为他们其中的一员吗？赶快抓紧机会 在国庆期间带上龙卡信用卡去境外享受一个不一样的假期吧。/ F5  . D9 a( G""  8 k1 s*  +  ' m* x- [& F$ ?- Q0  　　必备神器――龙卡全球支付信用卡$ T5 P& f. i: v% \$ @4 H( `; d$ W　　众多客户衷情的龙卡全球支付信用卡 到底有何魅力呢？且来看一下两笔境外消费的对比。如果在境外使用双币种信用卡消费1000英镑 这1000英镑将按照8月末英镑兑美元的汇率1.5442 折算为1544.2美元 再加上1.5%的兑换手续费 合计1567.36美元 计入双币种信用卡美元账户。还款时 按照6.4的汇率 则需要归还10031.10元人民币。但是 如果你选择的是龙卡全球支付信用卡 可免收外汇兑换手续费 直接按照英镑兑人民币的汇率9.8391 折算为9839.1人民币 足足节省了近200元。这样一计算 相信聪明的读者一定会做出明智的选择。. S! y) f; ]8 k3 x- D; L+ }+ t+ r/ A8 x- z; n8 v) Q1 O6 T　　优惠法宝――边游世界边赚钱. W* s  x  F| F. {0 d! q% M: E$ Z1 n* E9 W: ]　　没听错吧 境外消费或取现还能赚钱？如果你是龙卡信用卡客户 通过短信（CCHD#卡号后四位#010发送至95533）或“掌上龙卡”APP报名 就可以参加“龙卡信用卡玩转世界 境外消费或取现享6%返现奖励”活动。即日起至2016年6月30日期间每个自然月内 在境外消费/取现满6笔且每笔满等值600元人民币 即可获得当月境外消费/取现总金额6%的返现奖励（每持卡人每自然月最高奖励360元人民币）。6 P; O; W' ?. j5 D- a/ z1 B6 \% W9 b7 m% b. t* d  O　　如果你选择去日韩过节 则可使用龙卡JCB双币种卡或银联信用卡 在指定旅行社预订指定线路并出行 即可享受团费每单最高立减1000元优惠（每单2人起订）；如果使用龙卡日韩旅行信用卡（日本旅行卡JCB卡除外）每单可额外再减200元 更可在出行中畅享当地吃喝玩购海量特惠！: m: n8 V/ v! w""  ( ~  ^1 V; P7 p+ \4 C　　额度无忧――调额利器真便捷2 M$ V9 h$ s1 j% p* S9 z2 ]- Y| O0 o9 j& ?' u2 X' ?   　境外消费时额度不足怎么办？调额利器助您便捷申请提高临时额度 无忧消费。"" _1 ^% \( t3 k0 q7 O$ c1 c5 X"" A1 e# f. {/ K5 a1 P- E' }　　短信：通过在建行预留的手机号 编辑短信“CCTE#卡号后四位#申请额度”发送至95533申请临时额度调整。7 d  k$ Z2 t* ~"" k; {2 q- b4 ~: o) a8 G9 m) c/ Z　　网上银行：登录建行网上银行 依次点击“信用卡”―“信用卡额度调整”按提示完成即可。( O& W6 s& z* V+ N/ g- o+ ^2 R& V) v　　客服热线自助语音：拨打龙卡信用卡客服热线 根据语音提示依次输入“电话银行密码”―“需要调整的信用卡卡号后四位” 申请临时额度调整。; E) X7 D/ o& Z9 {; Z  @1 f. o贴心秘籍――微信“秘书”伴你行/ D| m   / E4 J' ]/ f6 m! x境外刷卡消费之时 如何能够时刻关注信用卡的“动态”呢？只需要关注“中国建设银行”微信银行 就能享受无“微”不至的龙卡信用卡服务。在微信银行绑定相应龙卡信用卡 即可实时收到境外刷卡的“外币消费/取现交易提醒” 交易时间、交易币种、交易金额、可用金额等一目了然点击“信用卡”板块 客户还可实时完成账单查询和还款、额度查询、积分查询、账单分期、约定账户设置、个人资料修改等九大功能操作。现在起信用卡绑定“中国建设银行”微信银行 即可参加信用卡达人指数测试 赢取信用卡账单免单机会；把活动分享到朋友圈 更可参与2888元年终大奖抽奖。6 J' v| s4 N* _7 m& D$ ~$ K' g"" j/ ^3 y. N: n建设银行| 信用卡| 出境旅游| 人民币| 手续费"|http://www.ngzb.com.cn/forum.php?mod=viewthread&tid=1244969&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline|2015-09-30
其他媒体|2038834380|zhidao_baidu|生活|ZHO|2015-09-30 22:28:01|东风悦达起亚k3车底有根管滴水是为什么|来自：手机知道汽车|http://zhidao.baidu.com/question/201536171159415005.html?fr=qlquick&entry=qb_list_default|2015-09-30
其他媒体|2038882620|zhidao_baidu|电子数码 > 手机/通讯-手机购买|ZHO|2015-09-30 22:59:02|东风悦达起亚k3空调排水管为什么排的那么慢|来自：手机知道汽车|http://zhidao.baidu.com/question/1820187860444069628.html?fr=qlquick&entry=qb_list_default|2015-09-30
其他媒体|2038934657|zhidao_baidu|游戏|ZHO|2015-09-30 23:33:02|起亚k3飞歌导航触屏没反应怎么处理|来自：手机知道汽车起亚k3飞歌导航触屏没反应怎么处理|http://zhidao.baidu.com/question/1670380398898474547.html?fr=qlquick&entry=qb_list_default|2015-09-30
其他媒体|2042509332|youku|生活|ZHO|2015-10-02 21:27:14|祝福祖国-生日快乐 重庆地铁员工串烧经典老歌|视频: 祝福祖国-生日快乐 重庆地铁员工串烧经典老歌|http://v.youku.com/v_show/id_XMTM0OTk3MDYyNA==.html|2015-10-02
其他媒体|2208192189|zhidao_baidu|文化/艺术|ZHO|2016-01-07 01:30:02|东风悦达起亚k3的平均油耗多少算正常|汽车|http://zhidao.baidu.com/question/1496898308189645379.html?fr=qlquick&entry=qb_list_default|2016-01-07
其他媒体|2208796233|zhidao_baidu|烦恼|ZHO|2016-01-07 11:23:02|东风悦达起亚k3汽车报价多少钱|汽车|http://zhidao.baidu.com/question/554620768218652412.html?fr=qlquick&entry=qb_list_default|2016-01-07
其他媒体|2208983235|bitauto|易车 > 问答 > 问题分类|ZHO|2016-01-07 13:10:02|东风悦达起亚k3的平均油耗多少算正常|东风悦达起亚k3的平均油耗多少算正常     提问者：易车网友 分类：  东风  买车  油耗  浏览[6]  2016-01-07 12:07  举报|http://ask.bitauto.com/detail/6068607/|2016-01-07
기타|2208988376|huanqiuauto|资讯 > 新闻|ZHO|2016-01-07 13:13:01|画面太美！ 2015年度最佳国民CP之汽车篇|2015年已挥手告别 年度最佳“国民CP”新鲜出炉 各种花式虐狗。星际有地球君与冥王星、政界有习大大与彭麻麻、娱乐圈有胡歌与霍建华……汽车圈有全新速锐与新帝豪。下面 我们一起来看看全新速锐/新帝豪这对家轿CP 到底谁更有魅力！		外形设计：均是年轻活力派  	       正如胡歌与霍建华这对CP 全新速锐与新帝豪虽已是业界前辈 但颜值丝毫不输鲜肉。前者前脸采用家族式“双飞翼”造型 搭配双幅镀铬条设计进气格栅、运动式前保险杠及LED日间行车灯等 辨识度颇高 再有双五辐造型铝合金轮毂、双边双出运动型尾排等时尚元素点缀 整车更是活力十足。后者在前脸、车身、尾部等细节均进行了优化 LED日间行车灯及后保险杠周边增加家族式回形纹 下进气栅格形状较现款更为隐蔽 镀铬条立体化等等 整车年轻不少。二者相遇 画面太美 叫人忍不住多看几眼。		装载能力：全新速锐略胜一筹	       中看还得中用。作为国民公认的实力派家轿 装载能力必须不俗。全新速锐拥有4680mm*1765mm*1490mm的长宽高、2660mm的轴距及450L的后备箱 直追B级车水平 多人出行也能舒适轻松 再搭配中央扶手箱、水杯卡位、手机盒等实用空间 实现物品随放随取 相当人性化。新帝豪长宽高为4631mm*1789mm*1470mm 轴距为2650mm 驾乘舒适感稍逊于全新速锐 不过也可以满足家庭的日常使用。		科技配置：全新速锐更显诚意	       在自主家轿市场 全新速锐与新帝豪这对搭档算是高科技、高逼格的典型。全新速锐素有“最安全自主轿车”之称 拥有ESP系统、内后视镜行车记录仪、TPMS胎压监测等几十项安全科技 同时搭载keyless系统、车载电视、10扬声器等多项智能配置 诚意十足。新帝豪则不及全新速锐到位 像CCS定速巡航、多媒体系统、全自动恒温空调等全新速锐标配科技 其只有中高配车型配备。下面 我们锁定两款车型的最高配展开比较 如下表：	 	    配置/车型    全新速锐1.5L自动旗舰型     2016款新帝豪1.3T CTV尊贵版      售价    9.59万    10.08万      PM2.5绿净系统    ●    —      360°全景影像    ●    —      发动机及空调遥控启闭    ●    —      Keyless智能钥匙    ●    ●      智能手表钥匙    ○    —      LED日间行车灯    ●    ●      ESP／ESC    ESP    ESC      TPMS胎压监测    ●    ●      主/副驾驶座安全气囊    主●/副●    主●/副●      前/后排侧气囊    前●/后—    前●/后—      前/后排头部气囊(气帘)    前●/后●    前●/后●      外后视镜电加热除霜    ●    ●      内/外后视镜自动防眩目    内○/外-    内-/外-      后视镜电动折叠    ●    —      行车记录仪    ○    ●      倒车雷达    6探头    4探头      GPS语音导航    ●    ●      车载数字电视    ●    —      车载蓝牙/电话    ●    ●      扬声器    10    6～7      CCS定速巡航    ●    ●      全皮型多功能方向盘    ●    ●      自动恒温空调    ●    ●      车内空气调节/花粉过滤    ●    —      G-Netlink3.0智能车载系统    ——    ●      CarPlay功能    ——    ●  		 	       可以看出 在配置方面全新速锐是比新帝豪要丰富 尤其是360°全景影像、PM2.5绿净系统、发动机遥控启闭等实用又时髦的科技 着实让全新速锐更占优势。就拿PM2.5绿净系统来说 通过过滤、吸附、净化三个步骤 轻松营造清新驾乘空间 拯救大家于雾霾深处。再看新帝豪 也就G-Netlink 3.0智能车载系统及CarPlay功能为整车平添了几分科技感。	       结语：从车本身来看 全新速锐比新帝豪更有吸引力 前者售价6.99万-9.59万 后者为6.98万-10.08万 同一价位区间 选择谁更实惠已无需多言。而且2016年1月1日——2016年1月31日期间 比亚迪还提供原本到2015年12月31日就结束的3000元惠民补贴 再加上购置税减半政策和比亚迪汽车金融公司“零等贷”活动 买辆全新速锐 省了好几千不说 月供还低 值得拥有！|http://www.huanqiuauto.com/news/20160107/849225_1.html|2016-01-07
其他媒体|2209213531|xcar_FORUM|论坛|ZHO|2016-01-07 15:29:01|一个老销售眼里的各种车评！|"之前写的一个评价车系感觉太繁琐 现在换个新的有评价 有美女图。大家要是有想咨询的车可以问我 帖子我就挑几个车型说说 不喜勿喷。丰田进口丰田耪ㄌ觳唤馐停盟溃业呐笥言谛薰淮考斯特之后对我说 妈的 怪不得温总理也用这玩意儿。广汽丰田的凯美瑞很棒 刹车没啥问题 价格公道质量也好 用不着批评。一汽的锐志和皇冠就不一样了 后刹车分泵时间长了活动的限位销子很容易锈蚀 直接后果就是“车到山前必有路 有路丰田刹不住”。v6缸水箱盖特别容易坏 不过也不算缺点 因为每一个漏防冻液的客户叫我来给他修车。我都是把他的水箱拆下来洗洗干净再装上去换个新盖子 收他一千多对他说“漏水了 我给你换个水箱。”变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后10％左右。福特。 进口福特没修过多少 房车修过但不多 钣金太差 拼缝和比亚迪一个水平。轮毂无一例外山寨感十足。合资福特 所谓的底盘和操控我没怎么感觉出来多厉害 和高尔夫差不多 做工钣金内饰水平一般 动力一般油耗偏高 经典福克斯节气门非常容易出问题 如果跑工地 电子节气门开度比例要不了多久就出问题 要换只有换总成 也就几千块 不贵但很烦 漏油情况不多 变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后30％左右。别克。 真别克 v6那种玩意儿 老车。油耗超高 漏油严重 气门饰盖和缸盖之间 也就是3缸与3缸两个夹脚没有垫子 只有打胶水 原车也是浇水 100多摄氏度老别克水箱风扇才会转 虽然我不知道是哪个煞笔设计到的这个温度 但是你可以想想 当水温到了100多度 那胶水能用多久？新别克 也就是大宇和欧宝换标车 漏油非常严重 洗了节气门就算不拆怠速也会上3000 仪器太差就无法匹配 仪器太好别人就要问你收钱 变速箱反应慢 降挡迟钝。变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后80％左右。日产日产是我这辈子见过最无语的车子 让人又爱又恨。你夸他内饰好吧 他外观差。你夸他动力强提速快吧他车子轻。你夸他油耗低吧他的机舱塑料用料小刀都能捅穿。你夸他配置高吧他大灯没透镜。你夸他隔音好吧他奶奶的每次抗日游行***暴动的时候 受伤最多的一定就是日产。不过有一个问题那就是 只要你开的是日产 开20年 都不会漏油漏水 除非你天天开出去撞 我真是服了他了 就是不漏！变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后0.005％左右。日产搭载的CVT变速箱很好 还有最重要是日产的发动机技术最成熟！斯巴鲁斯巴鲁这玩意好像只有进口的 除了brz之外都是全时四驱加水平对置发动机。曾经一款斯巴鲁力狮更是给我留下了“人车合一”的最好映像。缺点就是内饰穷 矮 丑。油漆硬度一般。打开发动机里面金属用料太差 这里点名斯巴鲁力狮水箱框架用两个手指头可以搬弯 这和吸能无关。离地间隙太小 车子特别容易托底碰石头 大灯没透镜看起来很难看。变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后20％左右 大多都是下面被石头刮漏的长城点名长城的哈佛H5是我这辈子见过质量最差的suv之一 轮胎很容易吃胎 什么球头橡胶罩子等小玩意儿更是不耐用 2.0na的发动机动力参数还不如奇瑞的1.6na 柴油皮卡车变速箱档把的皮套用的话顶多用个一年就掉色 车子停留久了打不着要一边打车一边就像做心脏起勃一样按它的手动油泵 很费劲儿。长城轿车大问题没啥 动力一般 低扭不足。由于哈佛h6销量太好 我也就不骂它了 我只是好奇1.5t没有直喷的增压算不算耍流氓？2d电影做成3d是不是也能骗过观众？点名某款老长城皮卡机油滤芯位置 发动机仓内朝上发动机后面 散热座子水管朝上 保养的时候没个半小时用三爪加公斤扳你拆不下来。介于长城不是越野就是跑工地 我评价已经很善良了 中国汽车吧的***不要喷我 变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后60％左右本田进口本田都是好车 很牛逼 但性价比不高。修的少就一代而过吧。国产本田 广汽的本田雅阁点名批评轮胎超级无敌特别非常容易轮胎扎钉漏气 不知道为什么 经常看见我徒弟补雅阁的胎 漏气就算了 还容易断轴 大灯没透镜太难看 车子金属材料一般 8代中控按键用得你手抽筋。东风的思域质量好 价格公道 底盘好 动力强 油耗低 缺点就是空调冷媒的橡胶管道容易出小洞 查漏怎么也查不出来 只有在特定角度漏气 妈的记得有一次全部拆下来在下面拼好放在水盆里打气都不漏 开出去没几天又漏了 我惹毛了 还了蒸发箱 压缩机和所有橡胶管道 ok 车主就从此以后再也不到我这里修车了。crv的刹车很线性 缺点暂时没发现 有的话就是太贵了。变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后10％左右。马自达进口马自达的车子很少出问题 来我这里都是做保险 就不说了。一汽马自达比如老马六 非常中庸 底盘不上不下 动力不上不下 油耗不上不下 外观不上不下 内饰不上不下 价格不上不下 空间不上不下 变速箱不上不下 名气不上不下 质量不上不下。 真他妈不上不下！不过有一点就是机盖支杆是在塑料水箱框架上 顶起来觉得不舒服 而且塑料水箱框架上装着水箱冷凝器 打灯 一撞换一大堆。长安马自达没遇到啥问题 都是来做保养 很丑性价比很低 就不说了 海南的搞过323不知道算不算马自达 车子的发动机气门顶筒要调节垫片 由于我技术太差 哪个人不幸地把自己的323给我绣的话无非两种情况。1:打不着 打着了怠速磨三天三夜不停的磨气门。 2:声音大 急加速吓得你尿都流到路腿上。变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后15％左右。大众这玩意儿我太有发言权了 进口大众好好使用97# 保养不差钱提前6/1周期做 机油用金美孚车子一般不会出问题。国产的老子特奶奶的现在就要开始骂人了 原谅我这里素质太低。卧槽上海大众 造10辆车就能在3年后漏10辆车 妈的上一趟高速后备箱里还要装上机油 轮胎什么牌子我就不铝耍1.6na发动机理机油口太小 保养没10分钟加不进去！加多了从油标尺抽油不出来！帕萨特b5 的bgc系列发动机三通管道真牛逼！造一个漏一个！换个新的开三个月又漏！换新的要蛮腰趴在机舱里照着电通换一个多小时 腰酸背疼还赚不到多少钱！减震非常容易漏油！一汽大众和上汽一样糟糕 就不多说了。高尔夫7代后悬挂简配 新速腾后悬挂简配！别的我就不隆Ｎ腋蠹医哺龉适拢乙话不崭缑嵌饰遥靶鄹纾陆荽锶绾危俊保宜怠耙孀泳吐蛉詹辽倏3年后不会漏油 大众一定会漏油的。”谁知道那***说:“漏油没关系 三年后说不定我就买新的了 大众车大气有面子。”我当时一听里怒了 对他说“你特么自己心里决定了还问老子干嘛！”。总结的说就是 大多数人买大众 钱多人傻价值观落后 请勿对号入座。变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后*******％左右。雪弗兰姨妈车质量还行 就是油耗高 动力差 车子安全性很好！大灯又他妈没什么透镜 低配没有esp 我无解了。进口姨妈的质量一般 油耗高 排量大 价格贵 na升功率一团糟 哪怕是8缸的雪弗兰也能被法拉利458的升功率爆出屎。合资姨妈点名科鲁兹内饰塑料感太强 光线采光不够 坐进去容易头晕 abs如果出问题了不解决一踩刹车就会熄火。漏油情况一般 变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后40％左右凯迪拉克作为为数不多的小众豪华品牌 凯迪拉克的性价比无疑是最高的。xts ats等等上搭载的高功率2.0T功率亮瞎！srx修过事故车 缺点就是配件问题 也可能是偶发问题但是一个地方反复发生各种问题 因为买的正厂配件 所以这种情况我个人不能接受。凯迪拉克没有什么显著缺点 变速箱的6at跟君威君越一个尿性 不过最近听说ats在金港跑过了进口328 感觉这些都无所谓 漏油不漏油没怎么注意看 因为修过的凯迪拉克都没有漏过。雷克萨斯雷克萨斯是我觉得就质量来说最好的车之一！还有一个就是奔驰！这两哥们的质量真的让人觉得狂拽霸帅酷耪ㄌ欤gs的发动机排量小 扭矩范围却能逆天！is动力、操控、外观、品牌独树一帜！ls质量稳定 隔音超一流！ct油耗低 价格低 维护保养贴心！lfa数量少 品质珍贵 跑圈必备！rx外观漂亮 内饰豪华！lx性价比虽然不高但是越野能力无出其右！总的来说 买雷克萨斯的人都是懂车的有钱人。不过介于这帖子是来黑车的 点名批评es系列油漆软！动力差！水箱盖很容易出问题！变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后0.0001％左右。雪铁龙雪铁龙的车子适合一个人开出去安安静静的兜风 人坐多了颠死人。我修过它的毕加索 觉得这车真的很渣 漏油漏水 关键是奇葩的水温表位置很容易让人看错 车内布局各种怪异 车子丑我就不说了 关键是售价还那么离谱。保养的时候找到空调滤芯 10个师傅就有5个找不到。点名批评雪铁龙世嘉发动机仓内排线混乱。而且变速箱技术落后还很费油 雪铁龙c5但是挺好 就是售价太离谱 而且毫无亮点。变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后80％左右。标致进口标志修过607 v6 通病没发现 也就是偶尔漏漏水 时常漏漏油。四个门拉手也就坏了三个 四个玻璃升降也就换了两个 别的也没啥 加点机油开一个月还剩一半而已。国产的东风标志除了车子丑 低配内饰差 变速箱渣 动力弱 油耗高 技术落后 配置低 外观丑之外也没有别的什么明显缺点。点名东风标志20 30 40 50漏油 漏水 漏空调冷媒 能漏的都漏 和大众3年漏光相比 如果大众3年新车10漏10 那么标致3年新车10漏9。变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后10086％左右。雷诺有人说雷诺就是日产 其实雷诺只是和日产有一些技术共享而已 和日产比技术还不行。雷诺的各种人机工程学设计近乎“反人类” 外观要么美得吓活人吓死 要么丑的把死人吓活。拉古娜古贝的四轮转向听着很牛逼其实开起来被奥迪35万那款高功率2.0t+夸托爆出屎 漏东西倒是不严重。牛逼轰轰的科雷傲性价比低不说还特么那么小=_= 不过梅甘纳系列还行！总的来说比psa的两个***车型好一点。变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后40％左右。奇瑞我大奇瑞总算出场了！别人都说奇瑞奇瑞 修车排队。其实都是放屁 不过这屁还是有一些道理的 为什么呢？因为奇瑞的发动机机构设计真的很得罪机修工 不挨骂活该！点名批评瑞虎 换个启动马达要拆进气歧管和水管等等等等 同样的工作要花别的车三倍的时间 全赚别人一样的钱 你说奇瑞挨不挨骂？新出的i auto平台的车型很棒！这里就不铝耍∑嫒鸬娜钡愦筇迨悄谑尾睿σ话悖侄渌傧涫指幸话悖忝榔嫒e5的内饰 两个字“好臭！” 漏油不多见但也有。变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后30％左右。帝豪全球鹰英伦其实他们都是一个品牌 除了ec7和ec8还行之外 其他的车都是渣。很多年以前我就说过 吉利的老板适合做生意不适合造车 旗下那么多品牌精品车型就那么两个 共同特点就是外观丑 动力差 装配工艺非常粗糙 牛逼吹的震天响 开起车来响震天！吉利的车质量还好！ec系列的销量和口碑都还行！点名批评吉利全球鹰gx7那神一样的动力和内饰 不多说了 说多了会吐。变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后20％左右。比亚迪比亚迪 我们先说优点吧 便宜 性价比高 早些年蓝天白云标的f3到处可见 比亚迪的车子优势在于“垂直整合” 很多零件都可以自己制造 便宜！所以性价比高得离谱！中国只有两个为中国人长脸的企业 一个叫华为 做手机的 一个叫比亚迪 造汽车的。缺点比亚迪也不少 外观差 内饰差 内饰用料就是凑个数 塑料拼缝不整齐 隔音不好 一脚刹车能把天窗绒板从后面滑到前面 小毛病多 品牌口碑烂 变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后30％左右。起亚起亚的车子真的是我见过用料差得车子中最突出的几个 看得见的地方增配 起亚使劲给你吹。看不见的地方减配 起亚使劲不让你黑。k2的面条轮胎有着无与伦比的垃圾质量 内饰烂 做工差 油漆没光泽 动力一般 变速箱马马虎虎。k3外形难看 大灯比概念车丑的多 黑色的后保险杠一脚能踢得掉下来 国外的朗动到国内变成k3后发动机还他么简配了……k4虽然不知道但一看名图觉得还不错 k5外观非常美丽就是不耐看 什么a柱异响 镜面轮毂高速跑断也时有发生。点名起亚智跑 如果你的车是智跑 做保养的时候叫师傅给你把车子顶起来 你看看他的悬挂 千万不要太伤心。变速箱、发动机、助力泵的油封、盖垫等等漏油几率新车三年后30％左右。奥迪：奥迪本不是什么豪华品牌 只不过在中国官车的成功挽救了奥迪 也让奥迪发现了在中国打高端牌的甜头 于是开始了高举高端的旗帜前进。奥迪最着名的招牌是发动机烧机油。这先天疾病来自大众。也在英国的评价中倒数第二 奥迪在三驾马车中无论是品位、品质、操控等都不占优 唯有主打科技感。奔驰：奔驰是汽车祖师爷 奔驰也用实际行动证明了 当汽车的祖宗决不能浪得虚名。无论碰撞测试还是各国分别进行的质量评估 奔驰都一直位居前列 绝不掉队。体现出了对汽车的真正理解真正实力。百年品牌 百年沉淀 实力不凡。当之无愧德系三驾马车之首。买奔驰任何一款车都不会有错 错的只是中外价格差别太大。不过沥青阻尼片、甲醛超标事件 给了奔驰下神坛的机会。宝马：三驾马车第二品牌 本来宝马在奔驰面前就是弱势 操控是弱势突围的手段 对操控观念的坚持也造就了宝马。宝马的质量控制并不如奔驰 在英国Autoexpress的发动机调查之中Mini荣登倒数行列之探花。宝马发动机功率不错 质量也只一般般 Autoexpress位列倒数第七。主打操控牌 让油耗低跟宝马交不了朋友。质量品质不如奔驰。以往各厂商都没有把客户的驾驶感受放在第一位 宝马的操控神主牌就高大地树立起来。现在操控优势已经不明显了。其实要论操控 高端操控跟宝马也没多大关系。要操控 所有轿车和SUV统统靠边|跑车上路。正好宝马就是生产轿车和SUV为主的。宝马Z是什么？Z3和奔驰SLK这种敞篷跑车都是马自达MX-5销售佳绩下刺激的产物。更何况宝马和公认最牛的WRC拉力赛的各个常务冠军车队搭不上边。宝马没那么神 一个以豪华为定位 以操控为卖点的家用车品牌。并不是说要把宝马贬低很普通合资车一样 宝马的操控和用料比普通合资车要强一些 但差距远没有价格那么大。保时捷：据说保时捷的品质很好 911很难驾驭。PANAMENA更像卖给装样子的暴发户的。这么贵的车 不易讨论。斯柯达：斯柯达是捷克和斯洛伐克的品牌 被大众收购之后 原有技术全部淘汰 就是大众的另一款孪生车。克莱斯勒：克莱斯勒被菲亚特收购了。克莱斯勒最著名的是JEEP。代表作是牧马人 不能用于实用的越野大玩具 当家用车来开的话 质量问题臭名远扬。这车是用来被车主折磨的 不是用来省心代步的。买这车需要明白这个道理。不图品牌不如看看北汽B40。便宜好多好多。菲亚特：意大利是超跑的故乡。家用车只有菲亚特。菲亚特是著名的“欧洲病车” 号称微车老大 但其产品在2012全世界汽车销量百强榜单之中 即使加上克莱斯勒的车型 也只有寥寥几辆。菲亚特比较小众 在国内的口碑还算不太好也不太坏 因为南京菲亚特时代 大家都没见过什么好车。菲亚特菲翔进入中国之后也出了断轴 还有发动机变速箱冒烟。同样配1.4T动力、DCT变速箱和扭力梁悬挂 比速腾便宜三万是有道理的。法拉利：法拉利虽然是菲亚特所属的投资集团旗下 但独立运营。有美国神车克尔维特C7在 昂贵的法拉利形象顿时贬值。法拉利林伯坚尼保时捷之类欧洲超跑都是坑有钱人的。原来不知道 后来再看性能对比标价就知道。参照物除了克尔维特还有路特斯（莲花）Elise。路虎 捷豹。卖给印度塔塔之后 在瓷器国反而身价暴涨 从优惠几万突然变成加价十几万。神！被列强抛来抛去的烫山芋在中国变成了香饽饽。阿斯顿马丁小马居然赖中国厂商生产的油门踏板是盗版材料 可笑的是中国生产的盗版材料配件居然6年以来没发生过任何故障 简直把阿斯顿马丁的脸打肿了。三菱：三菱在量产车上无论设计还是营销都很失败 但在基础工业上收获甚丰 不少国内外车企采购它的发动机配件 如发动机总成、涡轮增压器。和东南合作的V3菱悦卖了这么多年 机械搭配和操控精神上仍然让国产品牌10万以下A级车难以超越。三菱的机械不错 但卖货的本事却很低。三菱的缺点无非内饰粗糙点 毛病多点 价格稍贵点。其实安全、性能、油耗方面都不错 跟日产刚好相反。在傻子多的地方 骗钱都不会 那就没办法了。上汽之荣威和MG：外观设计无可挑剔 全系列车型国产车里面显得高端大气上档次。MG6和550开始及以上的车型底盘和用料值得称赞。虽然在英国评比中发动机倒数状元 但综合来讲在国内也是可靠的品牌 而且安全性是可靠的。但价格就不那么可靠了。上海人会营销 定价仅稍低于合资车 当合资车来卖 当然 比合资车来 还是厚道一些。特别是底盘 不输给主流合资同级产品 功力十足。550改款配DCT变速箱后降价 靠谱了很多 国产油老虎也变乖了不少。红旗国产第一品牌只有红旗一个能胜此任。红旗代表着中国国产车的最高技术和最高品质。红旗的任何一项水准直到目前为止仍比其他国产品牌高出一大班。拥有自主知识产权的6.0V12、4.0V8、3.0/2.5V6、2.0T、1.8T一系列高端发动机在孱弱的国产汽车工业中鹤立鸡群。丧心病狂的水军和无知的车盲黑白颠倒污蔑它们为丰田和大众发动机 实在可笑。没接触过H7的人容易带有色眼镜去看这俩车。即使有过接触的有些媒体人 依然喜欢带着有变形功能的有色眼镜 甚至主动担起颠倒是非的重任。实际上H7有不少挑战奥迪A6L的本钱。H7虽然无法撼动洋品牌C级车的地位 和国际高端品牌如奔驰宝马各方面都有潜在差距。但性价比绝对不低 车感不比奥迪A6L差。开红旗H7的气场比开同价位的宝马、奥迪还更威风煞气得多。奔腾如果不是一汽的管理层用行政思维代替市场经济来指导品牌运作 奔腾系列的销量远不是现在这般窝囊。主流级别的城市SUV之中 国产最佳技术最可靠仍然是X80 发动机变速箱底盘技术比其他国产SUV领先。贵有贵的道理。改款增加的1.8发动机B50值得一坑（十万买1.8改款马6还配后稳定杆 老马6改款后却阉割了） 今年的换代B70值得考虑。传说要增配2.0T的B90值得期待。得益于福特和马自达的技术 奔腾系列一直以来是品质和平衡性做得最优胜的国产车。不过反过来看 马自达上代技术开发的车型仍无其他国产品牌可以超越 唯有对国产车的发展再次抱憾。"|http://www.xcar.com.cn/bbs/viewthread.php?tid=25937507|2016-01-07
其他媒体|2223005067|webcars|降价信息|ZHO|2016-01-15 03:21:01|[郑州]  东风悦达起亚K5购车最高优惠现金3万元|"　　【万车网 郑州行情】近日 东风悦达起亚河南广发店内起亚K5最高优惠现金3万元 店内现车充足 颜色可选 欢迎试乘试驾 感兴趣的朋友不妨到店详询。详情优惠请见下表：　　近期火爆活动：　　【全城最低价 组团买新车】万车网团车活动火爆进行中（点击进入）　起亚K5郑州地区行情车型指导价（万元）现价（万元）优惠金额（万元）现车情况2016款 2.0T 自动PREMIUM23.9820.98↘3.00现车充足2016款 2.0T 自动LUXURY20.9817.98↘3.00现车充足2016款 2.0L 自动PREMIUM19.2816.28↘3.00现车充足2016款 2.0L 自动LUXURY17.5814.58↘3.00现车充足2016款 2.0L 自动GLS16.4813.48↘3.00现车充足2016款 2.0L 自动GL15.9812.98↘3.00现车充足2016款 1.6T 自动PREMIUM19.7816.78↘3.00现车充足2016款 1.6T 自动LUXURY18.0815.08↘3.00现车充足2016款 1.6T 自动GLS16.9813.98↘3.00现车充足2016年1月15日行情 车辆价格随时变动 敬请关注当地市场http://www.webcars.com.cn/zhengzhou/万车网制表您询问和购车时说明您是""万车网用户"" 会得到更好的服务！《点击可查看郑州地区东风悦达起亚4S店》　　2014款起亚新款K5在外观方面做了一些调整 其最大的变化集中在前脸细节方面 新车前大灯内部结构进行了调整 灯眉处增加了条形LED日间行车灯的设计 前脸的保险杠和新造型的雾灯边缘增加了镀铬装饰 同时下进气口的造型也进行了调整。而新增的2.0T车型 为了突出亮点 外观装饰有Turbo的标志 并且车尾处增加“TGDI”铭牌 展示涡轮增压车型的新身份。【2014款起亚K5 2.0T 外观】【2014款起亚K5 2.0T  外观】　　内饰设计方面 相较老款车型变化也不太大 中控台保留了向驾驶席倾斜角度的设计 采用了新样式的三辐方向盘 2.0T车型在内饰设计上也有别于普通车型 采用的是赛车式方向盘 底部为平直设计 为车内增加一些运动氛围。【2014款起亚K5 2.0T  内饰】【2014款起亚K5 2.0T 内饰】　　动力方面 新款K5新增2.0T涡轮增压车型 发动机最大输出功率为245马力 峰值扭矩达到350N·m 而普通的2.0L和2.4L车型动力系统则与老款相同。传动方面 除了2.0L入门级一款车型匹配手动变速箱之外 其余车型均使用了6速手自一体自动变速箱。　　经销商信息：　　经销商名称：河南普泽汽车销售服务有限公司　　经销商地址：河南郑州市郑东新区黄河南路和经北六路交叉口东北角　　经销商电话：****-******50|********　　声明：　　本文中涉及到的车型价格为万车网编辑在经销商处采集到的真实当日价格。由于汽车价格经常变化 并且为单一经销商的个体行为 所以价格仅供参考。具体价格请您致电或到店与经销商详细商谈。文中图片为车型实拍图 价格信息与图片拍摄地点无关。    本文导航         责任编辑：关鑫  关键词：起亚k5 k5报价及图片 k5怎么样 蒙迪欧 起亚k3 起亚k5怎么样 起亚k9 宾得k5 起亚k5最新报价 河南广发       查看车型   实时报价  参数配置  实拍图片  热点资讯  评分评论  万车知道"|http://www.webcars.com.cn/review/20160115/114114.html|2016-01-15
기타|2223634151|163_club|网易文化论坛-车迷闲聊|ZHO|2016-01-15 12:54:02|购买车辆时使用的什么类型的机油面。|雅鞍座套价格全包四季通用大众凌渡座套新迈腾座套高尔夫7专用座套新速腾新明锐坐套三防加厚版高尔夫7：淘宝价格680元；大众polo专用座套四季通用新polo 无级变速和自动挡哪个好汽车座套波罗车座套世嘉座套专用 苏格兰皮革+织物款：淘宝价格679元；全新福克斯座套经典福克斯两厢三厢汽车全包汽车专用四季夏季：淘宝价格510元；飞度卡罗拉威驰致炫XR-V缤智CR-V速腾骐达全包四季座套：淘宝价格519元；     独家真三防面料大众高尔夫6/新高尔夫7专用GTI苏格兰座套椅套：淘宝价格680元；全新福克斯座套经典福克斯两厢三厢汽车全包汽车专用四季夏季：淘宝价格359元；斯柯达明锐座套全包汽车专用坐套昕锐四季夏季冬季胜冰丝：淘宝价格509元；全包汽车坐套专用于大众新polo座套cross世嘉四季苏格兰：淘宝价格698元；     标致408专用汽车座套新桑塔纳新捷达坐套：淘宝价格465元；奥迪A3座套奥迪Q3座套奥迪A4L座套四季布艺全包专用座套：淘宝价格549元；丰田卡罗拉座套全包2014威驰致炫汽车坐套雷凌专用四季夏季：淘宝价格509元；雪铁龙世嘉座套全包三两厢汽车专用坐套四季CRV锋范：淘宝价格539元；     东风日产新阳光座套新轩逸全包座套夏季四季通用汽车坐套：淘宝价格952元；福特翼博座套全包翼搏汽车坐套新嘉年华专用三厢两厢福克斯：淘宝价格656元；奇瑞新qq座套骐达座套粉雅鞍凌派夏季仿皮雷凌夏季起亚k3座套新款：淘宝价格560元；新捷达专用汽车座套四季通用全包坐套桑塔纳朗逸专车定做：淘宝价格398元。小编结语不难发现这品牌的产品可以进行专属的制定 也有各种颜色的配制和选择。 途安机油的要求大众品牌的车辆很多都有他的专属机油 比如汽油发动机适用的型号有VW500、VW502、VW503、VW503.01、VW504 然而大排量的还需要参数HTHS≥3.5。主要起到的作用是节能、排气、清洁内部；柴油发动机使用的型号有VW505.00、VW505.01、VW506.00、VW506.01、VW507.00 主要针对于引擎设定。     途安机油的品牌     1、壳牌：主要选择的是灰壳的5W-40、 汽车之家二手车怎么样0W-40这两种型号的机油 由于灰壳的5W-30而大众品牌也可开始淘汰他。但是由于粘度比较低 所以用在新车里面的比较多。灰壳给我们带来的特点是噪音小、提高转速性能不好、提供动力性能不充分。      2、美孚1号：主要使用该品牌机油的型号有0W-40、5W-40 但是使用的都是金装美孚和金盖子美孚1号。虽然以前使用的0W-40、ESP5W-40这两种型号的机油比较多 由于这两款产生的噪音过大 提供动力不足地位也被其取代之。     3、嘉实多：主要也是使用的0W-40、5W-40这两种型号的机油 黑嘉5W-40这种型号虽然也在用 但是提供给车辆的保护系统是不很充分。由于该品牌的添加剂比较高端 因此提供的保护寿命也十分的长久。     4、福斯：使用最多的机油型号是泰坦超级合成5W-40 很多商家推荐说这款机油是非常适合大众车辆。因为该品牌在德国是专门为大众车辆提供润滑油产品的 在使用的过程中机油的消耗也非常合理。虽然提供的动力不如其他品牌 但是寿命和密封性却尤为的突出。     5、托库TR5、摩特8100X、300V、红线：这些被很多人称之为高价油 主要使用的型号也是5W-40。只要通过大众认证的40号产品 都可以在大众车上使用。这些高价油类型也有30号的使用 但是提供的耗油量很大。 途安机油的选择最初购买车辆时使用的什么类型的机油面 就可以继续的使用下去。如果你想换其他的机油试试 只要记住5W-40、0W-40这两种型号的机油 无论哪个品牌都有的 全车犀牛皮。大众品牌也是有自己专属的机油 为了爱车请慎重选择。小编结语通过对自己车辆的了解来进行机油的选择吧！|http://club.auto.163.com/bbs/auto_aaac/595206747.html|2016-01-15
其他媒体|2224025652|bitauto|易车 > 问答 > 问题分类|ZHO|2016-01-15 16:54:01|德系大众不考虑 韩系k3、和日系蓝鸟卡罗拉雷凌。哪个比较好！|德系大众不考虑 韩系k3、和日系蓝鸟卡罗拉雷凌。哪个比较好！     提问者：qcbjwx********  分类：  起亚  K3  买车  选车  浏览[6] 来自：易车手机客户端  2016-01-15 15:49  举报   德系大众不考虑 韩系k3、和日系蓝鸟卡罗拉雷凌。哪个比较好！求大神指教！|http://ask.bitauto.com/detail/6098654/|2016-01-15
其他媒体|2224653672|zhidao_baidu|电子数码 > 手机/通讯 > 通讯服务|ZHO|2016-01-15 23:43:02|怎样辨别东风悦达起亚k3是不是新车|生活常识|http://zhidao.baidu.com/question/1769300385850480380.html?fr=qlquick&entry=qb_list_default|2016-01-15
各大媒体|2256562316|bestb2b|全部信息|ZHO|2016-02-02 16:58:02|海兰德液压图混凝土车液压泵修理定州液压泵修理|"发布时间  2016年02月02日 国家地区   中国» 山东 » 济南    发布人 唐霞 公司  济南海兰德液压泵有限公司   地址  济南市历城区北园大街26号 网站  济南海兰德液压泵有限公司   邮件  ********@***.*** 手机  ***********   电话   ****-******36 QQ   **********    用户级别  普通会员       加入时间  2015年09月19日(距今136天)   精准匹配  混凝土车液压泵修理      报价  暂无报价     工程机械柱塞泵 柱塞泵马达 斜轴泵系列  德国力士乐A10VO| A4V| A11V柱塞泵系列 日本川崎 K3V| NV柱塞泵系列 日立系列：HPV116| HPV091国产CY14-1B柱塞泵等 泵在零件制造过程中 零件金属表面有一定的微观不平度(表面粗糙度)轴或孔存在的椭圆度与不直度 在金属表面发生初期相对运动时 泵零件间相对高速运动 此时摩擦副间会产生轻微的摩擦磨损 零件处于初期磨损阶段。 如果您对我们产品感兴趣 请拨打图片上面的电话 或者百度一下——海兰德液压泵客服电话联系我们 海兰德液压——您全程贴心的采购顾问 济南海兰德液压泵有限公司 公司主要经营液压泵、液压马达、液压测试仪、液压实验台的主要以液压泵（萨奥pv20系列）产品为主 其次还有川崎k3v系列、力士乐伊顿各系列产品及配件。公司成立十年来一直是在不断的学习引进国外的技术和经验。使我们的产品一直在不断地完善。越来越完美。 如果您对我们产品感兴趣 请拨打图片上面的电话 或者百度一下——海兰德液压泵客服电话联系我们 海兰德液压——您全程贴心的采购顾问 工程机械柱塞泵 柱塞泵马达 斜轴泵系列  德国力士乐A10VO| A4V| A11V柱塞泵系列 日本川崎 K3V| NV柱塞泵系列 日立系列：HPV116| HPV091国产CY14-1B柱塞泵等 泵在零件制造过程中 零件金属表面有一定的微观不平度(表面粗糙度)轴或孔存在的椭圆度与不直度 在金属表面发生初期相对运动时 泵零件间相对高速运动 此时摩擦副间会产生轻微的摩擦磨损 零件处于初期磨损阶段。 如果您对我们产品感兴趣 请拨打图片上面的电话 或者百度一下——海兰德液压泵客服电话联系我们 海兰德液压——您全程贴心的采购顾问联系我时请说明来自志趣网 谢谢!"|http://www.bestb2b.com/business_91824962.htm|2016-02-02
其他媒体|2267204859|zhidao_baidu|游戏|ZHO|2016-02-09 00:47:12|起亚k3gls和比亚迪速悦那个好|汽车|http://zhidao.baidu.com/question/393978317616871405.html?fr=qlquick&entry=qb_list_default|2016-02-09
其他社区|2267889001|360wenda|待解决问题|ZHO|2016-02-09 14:35:01|英朗.卡罗拉.k3.哪个比较好.18岁开|英朗.卡罗拉.k3.哪个比较好.18岁开Ooo苏陌ooO10级分类： 汽车被浏览38次4分钟前请微博专家回答检举|http://wenda.haosou.com/q/1454995786494167|2016-02-09
其他媒体|2268564655|mobile01|新進文章|ZHO|2016-02-09 23:31:01|LEXUS ct200h&is200t 的一些疑問|各位前輩好小弟現在開的是ford focus mk3  因為努力工作也存了一筆錢 準備要換新車了從 BENZ gla180  BMW X1 福斯sportsvan  一直看到lexus ct200h 和is200t想請問目前 lexus折價高嗎？ 大概都是定價折多少呢？？ 另外ct200h 菁英款本身配備足夠嗎？因為本人工作關係 很常全台灣各地跑 市區也很常跑  所以主要是看上ct200h的省油性本人不習慣飆車 高速公路開車也常在 110~120左右 偶爾超車 也會跑山路 不知道ct200h是否有力 不用快只要不要爬不上坡就好！看他的相關報導有sport模式 不知道菁英版也有嗎？後座部分也有聽朋友說非常的小 很不推薦 但目前只有我跟我女友使用 後座部分不常載人 我預計170~175左右的人能坐就好 在高的自己去想辦法ＸＤ  想詢問是真的非常的不夠嗎？ 小弟本身也是175另外他屬於油電車款 不知道會不會常有些零件壞掉呢？ 另外又看到us200t是覺的外型十分帥氣 所以也一起加進了比較清單再來lexus的保養部分 不知道會不會很貴？ 還有零件更換會不會也很昂貴呢？再麻煩有購買lexus車款的前輩們可以分享一些建議了！ 非常感謝另外如果有推薦業務也可以一起推薦給我喔！！|http://www.mobile01.com/topicdetail.php?f=346&t=4704852|2016-02-09
各大媒体|2278298514|enorth|汽车频道|ZHO|2016-02-15 16:30:02|悦达起亚k3现车优惠4万 k3全系折扣巨惠|悦达起亚k3现车优惠4万 k3全系折扣巨惠 来源：网上车市　作者：　2016-02-15 13:52:19　编辑：杨辰    　　【网上车市天津滨海行情.原创】近日获悉 东风悦达起亚k3现车到店 东风悦达起亚k3最新促销价格全系优惠4万。东风悦达起亚k3配置丰富手续齐全 具体颜色和配置请致电商家咨询 更多优惠尽在北京万仁众泰汽车销售有限公司 如您对本车感兴趣 欢迎致电咨询 购车热线：　　*********** 刘经理　　具体车型以及价格如下：　　本车报价：　　外观方面 东风悦达起亚k3在前脸的设计上十分突出力量感和线条的精炼 采用起亚旗舰车型K9的镀铬直瀑式竖条进气格栅 视觉感受更为大气、稳健 后尾组合尾灯和外后视镜集成转向灯都采用LED设计 再配合LED日间行车灯 彰显出浓厚的科技感以及时代感。　　细节方面 东风悦达起亚k3的超长轴距更打造出同级别最大乘用空间 充分保障了驾乘舒适性。K3还配备了电动通风真皮座椅、双区恒温空调、一键启动、高级音响系统等同级罕见的科技 充分体现出K3配置的丰富和越级。　　内饰方面 东风悦达起亚K3简约内饰 完满组合时尚先锋梦之队。K3内饰做工精致 真皮座椅、方向盘、门护板、仪表盘等皮质包裹 触感细腻高贵 工艺超越同级。K3的配置套餐也极具智能感 与K3族群“科技控”的前瞻审美观无缝衔接。　　配置方面 东风悦达起亚k3还搭载了起亚最新的1.6L伽马D-CVVT和1.8L Nu D-CVVT两款发动机 最大功率分别达到128马力和146马力 动力强劲且燃油经济性突出。配合先进的6速手自一体变速箱 操控随心 能很好的开发车主驾驭热情。【网上车市天津滨海行情.原创】　　更多详情请点击： http://binhai.cheshi.com/ 网上车市滨海车市 　　温馨提示：以上 购车 优惠信息由天津滨海综合 经销商 提供 仅供 购车 参考；由于行情因素价格浮动较大 具体车辆成交价格请致电商家获取最新报价；优惠行情可查阅网上车市天津滨海 经销商 报价后台 告知对方信息来源于网上车市将有更多优惠。|http://auto.enorth.com.cn/system/2016/02/15/030808335.shtml|2016-02-15
其他媒体|2278944842|bitauto|易车 > 问答 > 问题分类|ZHO|2016-02-15 22:50:02|起亚k4报价东风悦达起亚k3怎么样|起亚k4报价东风悦达起亚k3怎么样     提问者：易车网友 分类：  起亚  K4  买车  报价  浏览[6]  2016-02-15 21:46  举报|http://ask.bitauto.com/detail/6195246/|2016-02-15
其他媒体|2298528958|zhidao_baidu|烦恼|ZHO|2016-02-26 00:41:02|长安欧诺2o16a2k3报价?|汽车|http://zhidao.baidu.com/question/1693279502682001308.html?fr=qlquick&entry=qb_list_default|2016-02-26
其他媒体|2298782319|zhidao_baidu|电脑/网络 > 电脑装机|ZHO|2016-02-26 05:05:01|东风悦达起亚k3在110码的时候急转弯会不会翻车…|汽车|http://zhidao.baidu.com/question/1821151317874986708.html?fr=qlquick&entry=qb_list_default|2016-02-26
其他媒体|2299496082|bitauto|易车 > 问答 > 问题分类|ZHO|2016-02-26 14:29:01|东风悦达起亚k3在110码的时候急转弯会不会翻车…|东风悦达起亚k3在110码的时候急转弯会不会翻车…     提问者：易车网友 分类：  东风  其他  浏览[6]  2016-02-26 13:25  举报|http://ask.bitauto.com/detail/6233100/|2016-02-26
其他媒体|2299951586|bitauto|汽车行情 RSS|ZHO|2016-02-26 18:48:01|娇小干练、舒适性高 爱你没商量的小2|"品牌：  起亚  车款：  起亚K2三厢 1.4L 自动 GLS  油耗：8.1L 评分：       外观   内饰   空间   动力   操控   配置   性价比   舒适度                油耗：今天刚加的油 到月底还有好几天 2月份全月大概油耗在每公里0.45元 每月大概跑600公里左右 总体花费在350-400元之间 总体来说还是较为省油的 最近因为天气越来越暖和 所以油耗下降很多 而且春节期间跑的也多些。    外观：外观我想是很多车友选k2首选的 我也是外观控 对于k2的前脸特别喜欢 虽然车身流线型与k3|k4相比较差了很多 但整体不失比例 无论哪个角度来看 都没有不协调感。轮毂不是镜面的 但我认为也不差 而且全铝的。    内饰：内饰的塑料感还是明显的 而且到现在我的车子里面 还是有一点气味 所以每次开车前会开窗通气 因内饰是全黑的 所以容易脏 经常性的打理 用手摸上去 塑料感不是特明显。  空间：整体空间 驾驶和副驾驶空间还是蛮大的 可能是我向后放倒的原故 后排三座空间可以 就是腿放下后空间不是很舒服 需要斜着放 时间长了有点酸 但座位不小 坐上去后不显的小 后备箱还是较大的 我里面放了很多的东西 主要还是常备的工具和一些物品 过年送节放礼品 几家的一起放里 都不显的挤。  动力：对于小2的动力 我认为还是不错的 1.4的排量 不要指望它能给你带来多大的惊喜 主要还是起步有点肉肉的 不会给予太强的动力 其实舍的给油 但我认为没有必要 缓慢起步 也是安全行车的一部分。  操控：用了两年了 单手都可以随意操控 但出于安全 还是双手 说明方向盘还是较轻的 但底盘还是有点轻 在40码拐弯时还是有点飘的感觉 不过在高速上 均速提速后 车子整体还是很科稳的 就是噪音大了些 有些受不了 不过习惯就好了。  配置：我自己这款配置不是很多 基本常用都有 CD用的不多 主要还是听广播的多 没有导航 也不喜欢加那个东西 感觉实在的还是倒车雷达 后视窗加热功能。  性价比：车子用了快两年了 基本已经适应了自己车子的各项性能 基本够用 对于一些特殊的功能 我自己给加配上去 以实用为主 当时在选小2前 还是作了功课的 当时看重速锐、飞度 但后来都没有选中 主要还是喜欢小2的外观和实用性。  舒适度：舒适度一般化了 毕竟不是真皮座椅 是针织座椅 而且后排座位不能调节 长时间坐有些不舒服感 计划今年有钱的话 想换套真皮座椅 提高一些档次的同时 也让车子的舒适度提升一下。  当前里程：13900 公里   裸车价：800400万   芜湖  2014年4月购车  经销商： 芜湖顺易起亚        k2买回来快2年了 跑的公里数不多 但总体来说没有掉链子过 对于自己当初的选择还是满意的 时尚的外观 自动挡车型配备挡位提示功能 价格便宜 在同级别的紧凑型车型来说都是性价比最高的。某宝上买的座垫 质量不是很好 先凑合着用吧。来张侧面照加油前跑的公里数CD有点不上档次 但还是较为实用性的。    车主过往口碑  购车1年我的小2 我自豪    0"|http://bitauto.feedsportal.com/c/33450/f/584188/s/4dde2b7b/sc/17/l/0Lbaa0Bbitauto0N0Ck20Cthread0E87481410Bhtml/story01.htm|2016-02-26
기타|2402771582|Autohome review|혼다 어코드(雅阁)|ZHO|2016-04-24 00:35:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=67&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-04-24
其他媒体|2402815777|youku|汽车|ZHO|2016-04-24 01:11:01|颜值爆表 2017款丰田卡罗拉50周年版||http://v.youku.com/v_show/id_XMTU0NTYwMzk3Mg==.html|2016-04-24
기타|2402915236|Autohome review|혼다 어코드(雅阁)|ZHO|2016-04-24 02:49:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=68&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-04-24
기타|2403346613|Autohome review|혼다 어코드(雅阁)|ZHO|2016-04-24 12:20:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=69&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-04-24
기타|2403422926|Autohome review|혼다 어코드(雅阁)|ZHO|2016-04-24 13:23:02|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=70&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-04-24
기타|2410452882|Autohome review|혼다 어코드(雅阁)|ZHO|2016-04-28 00:18:14|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=100&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-04-28
기타|2411324048|Autohome review|혼다 어코드(雅阁)|ZHO|2016-04-28 12:46:06|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=101&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-04-28
其他媒体|2411423996|bitauto|易车 > 问答 > 问题分类|ZHO|2016-04-28 13:49:01|比亚迪“宋”怎么样？油耗高吗？手动低配的十万内能搞定吗？有...|比亚迪“宋”怎么样？油耗高吗？手动低配的十万内能搞定吗？有没     提问者：YCAPP*******RJW2  分类：  起亚  K3  买车  车型  浏览[2] 来自：易车手机客户端  2016-04-28 12:36  举报   比亚迪“宋”怎么样？油耗高吗？手动低配的十万内能搞定吗？有没有车主啊 说说下感觉怎样？不行的话只能买k3了|http://ask.bitauto.com/detail/6488355/|2016-04-28
기타|2412005946|Autohome review|혼다 어코드(雅阁)|ZHO|2016-04-28 18:58:03|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=104&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-04-28
其他媒体|2412102689|bitauto|易车 > 问答 > 问题分类|ZHO|2016-04-28 19:53:04|k3 自动 gls 哈弗h6自动精英版  选哪|k3 自动 gls 哈弗h6自动精英版  选哪     提问者：熊旭  分类：  起亚  K3  买车  选车  浏览[2] 来自：汽车报价大全  2016-04-28 18:48  举报   相关车型：起亚K3|http://ask.bitauto.com/detail/6489854/|2016-04-28
기타|2412213157|Autohome review|혼다 어코드(雅阁)|ZHO|2016-04-28 20:57:05|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=103&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-04-28
기타|2476115533|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 00:16:27|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=177&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-06-02
기타|2476125700|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-02 00:22:05|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=140&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-06-02
기타|2476143189|Autohome_review|랑동(朗动)|ZHO|2016-06-02 00:32:01|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=213&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-06-02
기타|2476145149|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 00:33:02|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=121&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-06-02
기타|2476145176|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 00:33:02|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=103&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-06-02
기타|2476145180|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 00:33:02|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=100&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-06-02
기타|2476163904|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 00:45:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=118&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-06-02
기타|2476187494|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 01:00:04|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=203&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-06-02
기타|2476187686|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 01:00:04|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=7&piap=0 2886 0 0 2 0 0 0 0 0 1#20151015|2016-06-02
기타|2476213031|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-02 01:17:05|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=141&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-06-02
기타|2476217617|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-02 01:21:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=214&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-06-02
기타|2476217722|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-02 01:21:01|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=170&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-06-02
기타|2476226488|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 01:27:33|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=123&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-06-02
기타|2476226537|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 01:27:33|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=105&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-06-02
기타|2476226544|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 01:27:33|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=102&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-06-02
기타|2476262574|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 01:54:02|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=204&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-06-02
기타|2476262765|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 01:54:02|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=9&piap=0 2886 0 0 2 0 0 0 0 0 1#20151015|2016-06-02
기타|2476306162|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 02:34:01|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=119&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-06-02
기타|2476330500|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 03:00:02|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=178&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-06-02
기타|2476535891|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 07:47:09|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=179&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-06-02
其他媒体|2476558216|bitauto|易车 > 问答 > 问题分类|ZHO|2016-06-02 08:11:03|11万到十二万从各种角度来看 哪种紧凑型车好！ 就现代|11万到十二万从各种角度来看 哪种紧凑型车好！ 就现代     提问者：点击查看更多！  分类：  买车  选车  浏览[0] 来自：汽车报价大全  2016-06-02 07:10  举报   11万到十二万从各种角度来看 哪种紧凑型车好！ 就现代朗动1.6L手动尊贵型 和领动1.6手动致炫活力型 和k3手动高配 从空间实用 外观 安全 油耗 综合考虑 买哪个好 |http://ask.bitauto.com/detail/6616884/?leads_source=p029001|2016-06-02
기타|2476563115|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 08:15:01|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=120&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-06-02
기타|2476596707|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-02 08:46:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=215&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-06-02
기타|2476596813|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-02 08:46:02|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=171&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-06-02
기타|2476730464|Autohome_review|뉴 보라(宝来)|ZHO|2016-06-02 10:18:03|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=182&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-06-02
기타|2476750820|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 10:30:01|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=180&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-06-02
기타|2476785720|Autohome_review|랑동(朗动)|ZHO|2016-06-02 10:51:02|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=215&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-06-02
기타|2476801231|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 10:59:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=121&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-06-02
기타|2476808638|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-02 11:04:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=216&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-06-02
기타|2476808773|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-02 11:04:02|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=172&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-06-02
기타|2476859600|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 11:32:02|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=122&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-06-02
기타|2476859640|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 11:32:02|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=104&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-06-02
기타|2476859643|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 11:32:02|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=101&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-06-02
기타|2476859728|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 11:32:02|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=8&piap=0 2886 0 0 2 0 0 0 0 0 1#20151015|2016-06-02
기타|2476898207|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-02 11:53:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=142&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-06-02
기타|2476914509|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 12:02:01|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=181&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-06-02
기타|2476914576|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 12:02:01|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=122&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-06-02
기타|2476938366|Autohome_review|뉴 보라(宝来)|ZHO|2016-06-02 12:15:01|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=183&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-06-02
기타|2476941370|Autohome_review|랑동(朗动)|ZHO|2016-06-02 12:16:52|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=216&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-06-02
기타|2477028753|Autohome_review|랑동(朗动)|ZHO|2016-06-02 13:12:02|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=217&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-06-02
기타|2477052877|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-02 13:28:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=217&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-06-02
기타|2477052922|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-02 13:28:02|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=173&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-06-02
기타|2477149043|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 14:29:01|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=205&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-06-02
기타|2477149143|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 14:29:01|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=124&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-06-02
기타|2477149171|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 14:29:01|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=106&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-06-02
기타|2477192233|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 14:55:02|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=103&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-06-02
기타|2477192566|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 14:55:02|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=10&piap=0 2886 0 0 2 0 0 0 0 0 1#20151015|2016-06-02
기타|2477216968|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-02 15:11:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=143&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-06-02
기타|2477274853|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 15:45:02|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=182&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-06-02
기타|2477274912|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 15:45:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=123&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-06-02
기타|2477432099|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 17:13:02|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=183&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-06-02
기타|2477486345|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-02 17:42:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=219&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-06-02
기타|2477486439|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-02 17:42:02|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=174&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-06-02
기타|2477488782|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 17:43:01|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=207&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-06-02
기타|2477488875|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 17:43:01|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=126&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-06-02
기타|2477488917|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 17:43:01|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=108&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-06-02
기타|2477488924|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 17:43:01|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=105&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-06-02
기타|2477497541|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 17:47:32|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=124&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-06-02
기타|2477529604|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 18:04:01|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=12&piap=0 2886 0 0 2 0 0 0 0 0 1#20151015|2016-06-02
기타|2477664493|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-02 19:19:01|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=175&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-06-02
기타|2477680483|Autohome_review|뉴 보라(宝来)|ZHO|2016-06-02 19:28:02|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=184&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-06-02
기타|2477685713|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 19:32:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=125&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-06-02
기타|2477730664|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 20:00:01|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=185&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-06-02
기타|2477777787|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-02 20:30:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=126&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-06-02
기타|2477984838|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 22:33:01|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=208&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-06-02
기타|2477985236|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 22:33:02|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=127&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-06-02
기타|2477985363|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 22:33:02|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=109&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-06-02
기타|2477985387|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 22:33:02|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=106&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-06-02
기타|2478002340|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-02 22:43:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=144&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-06-02
기타|2478029811|Autohome_review|K3(起亚K3)|ZHO|2016-06-02 22:59:01|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=13&piap=0 2886 0 0 2 0 0 0 0 0 1#20151015|2016-06-02
기타|2478121340|Autohome_review|아반떼 AD(领动)|ZHO|2016-06-02 23:57:03|2016年06月02日 发表了口碑|来自：手机汽车之家  2016年06月02日 发表了口碑  口碑   《外观拉风 配置足够 整体性价比还是不错的。》           【最满意的一点】外观很拉风 现在路上还很少见 大轮毂。日间行车灯很高大上 自动头灯也很高端。中控台是软的 车内显示屏清晰度很高。倒车影像有随动辅助导线。很方便。车内音响很赞 我喜欢听音乐 完全满足我的要求。【最不满意的一点】后排不能放倒 这个真心很郁闷 这个放倒真的很难吗？这几天B柱内有异响 这还是新车呀 哎。。过几天去4s看看 希望不是啥大问题。另外胎噪确实大 我想跟轮胎大也有关系吧。悬挂还是有点硬 不过在接受范围内。【空间】空间同级别还是有优势的 中间无凸起。【动力】动力够用 现在用的eco模式【操控】转向精准 没啥虚位。【油耗】表显6 肯定是不准的 等下次油表亮再算算。【舒适性】还可以 家用够了。【外观】满意【内饰】做工还是比较好的 接缝均匀。【性价比】性价比高【为什么最终选择这款车？】同级别都看了 也试驾了 福克斯空间太小 科鲁兹都说油耗高 新英朗有点老气 卡罗拉没esp 思域根本没现车 看来看去家用也就韩系车了。【其他描述】换车的想法去年就有了 但是一直没有付诸行动 一是因为暂时有车开 二是今年上市新车多 想再等等 经常看论坛 心里已经有了几个备选 英朗 老表刚买的 开始觉得性价比很高 后来发现新旧差别很大 就pass了。福克斯外观不错 但是同事有好几辆 不想买一样的。k3性价比很高 优惠很大 但是新款感觉你没老款好看。看到最后就是领动了 配置高 外观拉风 总体性价比很高。|http://k.autohome.com.cn/spec/25701/view_1148059_1.html?st=1&piap=0 3959 0 0 2 0 0 0 0 0 1#20160602|2016-06-02
기타|2497827395|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-14 00:28:18|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=15&piap=0 982 0 0 2 0 0 0 0 0 1#20160612|2016-06-14
기타|2497836019|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 00:31:01|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=167&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-06-14
기타|2497836076|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 00:31:01|2016年05月19日 发表了质量评价|2016年05月19日 发表了质量评价  质量   【行驶过程】  刹车时有异响-车辆前部  【内饰】  随车脚垫会滑动或污损       来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=149&piap=0 2886 0 0 2 0 0 0 0 0 1#20160519|2016-06-14
기타|2497836087|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 00:31:01|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=146&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-06-14
기타|2497836359|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 00:31:02|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=55&piap=0 2886 0 0 2 0 0 0 0 0 1#20151015|2016-06-14
기타|2497871283|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-14 00:55:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=193&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-06-14
기타|2497890991|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 01:07:24|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=170&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-06-14
기타|2497891033|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 01:07:24|2016年05月19日 发表了质量评价|2016年05月19日 发表了质量评价  质量   【行驶过程】  刹车时有异响-车辆前部  【内饰】  随车脚垫会滑动或污损       来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=152&piap=0 2886 0 0 2 0 0 0 0 0 1#20160519|2016-06-14
기타|2497891036|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 01:07:24|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=149&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-06-14
기타|2497891176|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 01:07:30|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=57&piap=0 2886 0 0 2 0 0 0 0 0 1#20151015|2016-06-14
기타|2497891206|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 01:07:31|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=43&piap=0 2886 0 0 2 0 0 0 0 0 1#20160604|2016-06-14
기타|2497891271|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 01:07:31|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=20&piap=0 2886 0 0 2 0 0 0 0 0 1#20160608|2016-06-14
기타|2497934144|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 01:38:03|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=58&piap=0 2886 0 0 2 0 0 0 0 0 1#20151015|2016-06-14
기타|2497934175|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 01:38:03|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=44&piap=0 2886 0 0 2 0 0 0 0 0 1#20160604|2016-06-14
기타|2497934250|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 01:38:03|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=21&piap=0 2886 0 0 2 0 0 0 0 0 1#20160608|2016-06-14
기타|2497935313|Autohome_review|BYD S6(比亚迪S6)|ZHO|2016-06-14 01:39:01|2016年04月01日 发表了口碑|来自：汽车之家iPhone版  2016年04月01日 发表了口碑  口碑    《空间大就不用说了 没有之前担心的动力不足 感觉动力够用》           【最满意的一点】空间 配置 虽然2.0手豪（不想要天窗 应人而异）但是后期选装自装也是感觉很霸气 好多十多万的车都没有的配置  心里美滋滋～【最不满意的一点】目前就发现右后轮起步有点异响 但是说来也怪  每次到4s店就没有了 去了四五次都不响了 回家没几天又继续  好邪～【空间】前几天去了东北  （有贴） 后面气垫床谁俩人（178cm）没问题  还能装点东西～【动力】没有网上说的那么肉  我只想说只要舍得给油什么车都不肉【操控】开的还不错  就是刚开始开离合太高不习惯  现在习惯了 感觉很透  油门也挺灵活  （之前在部队开猛士） 开小六感觉 很棒【油耗】比预计要低可能跑长途的 以前市区差不多9个油还能接受 这次高速回来平均降到8.7 不管多少2.0这么大的车 只要不超十个油都能接受【舒适性】椅子倍舒服 以前猛士没法比  也不能比 不是一个级别 感觉比朋友的k3舒服多了！【外观】外观挺不错的  不过现在出来好的新车自然小六要逊色不少  不过自己折腾加装踏板 牛头杠 行李架 （准备换Q5大灯和仿宝马LED尾灯）【内饰】内饰除了座椅和方向盘很满意 其他都很一般般吧！【性价比】性价比就不说了直接满分  这么大的车裸车7w多块钱 去哪找？【为什么最终选择这款车？】其实购车前一直看中h6  但是资金有限（不想贷款）全身就10w  后来看了好多款  家里差点让买了宝骏560  和陆丰x7（家里支持资金）但是最后还是选择了s6 因为家里不喜欢比亚迪 这个名字（大家好多都懂的）说十几万宁愿买个CRV  不过我不喜欢日产（还是应人而异）【其他描述】|http://k.autohome.com.cn/spec/18563/view_1041472_1.html?st=184&piap=0 2088 0 0 2 0 0 0 0 0 1#20160401|2016-06-14
기타|2497971536|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 02:09:01|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=171&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-06-14
기타|2497971574|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 02:09:01|2016年05月19日 发表了质量评价|2016年05月19日 发表了质量评价  质量   【行驶过程】  刹车时有异响-车辆前部  【内饰】  随车脚垫会滑动或污损       来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=153&piap=0 2886 0 0 2 0 0 0 0 0 1#20160519|2016-06-14
기타|2497971580|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 02:09:01|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=150&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-06-14
기타|2497971974|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 02:09:02|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=59&piap=0 2886 0 0 2 0 0 0 0 0 1#20151015|2016-06-14
기타|2498001911|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 02:36:02|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=45&piap=0 2886 0 0 2 0 0 0 0 0 1#20160604|2016-06-14
기타|2498001963|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 02:36:02|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=22&piap=0 2886 0 0 2 0 0 0 0 0 1#20160608|2016-06-14
기타|2498237975|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 07:44:01|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=172&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-06-14
기타|2498238031|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 07:44:01|2016年05月19日 发表了质量评价|2016年05月19日 发表了质量评价  质量   【行驶过程】  刹车时有异响-车辆前部  【内饰】  随车脚垫会滑动或污损       来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=154&piap=0 2886 0 0 2 0 0 0 0 0 1#20160519|2016-06-14
기타|2498238039|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 07:44:01|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=151&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-06-14
기타|2498284592|Autohome_review|뉴 보라(宝来)|ZHO|2016-06-14 08:32:01|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=219&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-06-14
기타|2498290476|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 08:37:02|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=173&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-06-14
기타|2498290513|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 08:37:02|2016年05月19日 发表了质量评价|2016年05月19日 发表了质量评价  质量   【行驶过程】  刹车时有异响-车辆前部  【内饰】  随车脚垫会滑动或污损       来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=155&piap=0 2886 0 0 2 0 0 0 0 0 1#20160519|2016-06-14
기타|2498290516|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 08:37:02|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=152&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-06-14
기타|2498290869|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 08:37:03|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=61&piap=0 2886 0 0 2 0 0 0 0 0 1#20151015|2016-06-14
기타|2498290910|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 08:37:03|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=47&piap=0 2886 0 0 2 0 0 0 0 0 1#20160604|2016-06-14
기타|2498290947|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 08:37:03|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=24&piap=0 2886 0 0 2 0 0 0 0 0 1#20160608|2016-06-14
기타|2498371173|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-14 09:41:04|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=16&piap=0 982 0 0 2 0 0 0 0 0 1#20160612|2016-06-14
기타|2498376632|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-14 09:45:01|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=194&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-06-14
기타|2498383836|Autohome_review|BYD S6(比亚迪S6)|ZHO|2016-06-14 09:49:02|2016年04月01日 发表了口碑|来自：汽车之家iPhone版  2016年04月01日 发表了口碑  口碑    《空间大就不用说了 没有之前担心的动力不足 感觉动力够用》           【最满意的一点】空间 配置 虽然2.0手豪（不想要天窗 应人而异）但是后期选装自装也是感觉很霸气 好多十多万的车都没有的配置  心里美滋滋～【最不满意的一点】目前就发现右后轮起步有点异响 但是说来也怪  每次到4s店就没有了 去了四五次都不响了 回家没几天又继续  好邪～【空间】前几天去了东北  （有贴） 后面气垫床谁俩人（178cm）没问题  还能装点东西～【动力】没有网上说的那么肉  我只想说只要舍得给油什么车都不肉【操控】开的还不错  就是刚开始开离合太高不习惯  现在习惯了 感觉很透  油门也挺灵活  （之前在部队开猛士） 开小六感觉 很棒【油耗】比预计要低可能跑长途的 以前市区差不多9个油还能接受 这次高速回来平均降到8.7 不管多少2.0这么大的车 只要不超十个油都能接受【舒适性】椅子倍舒服 以前猛士没法比  也不能比 不是一个级别 感觉比朋友的k3舒服多了！【外观】外观挺不错的  不过现在出来好的新车自然小六要逊色不少  不过自己折腾加装踏板 牛头杠 行李架 （准备换Q5大灯和仿宝马LED尾灯）【内饰】内饰除了座椅和方向盘很满意 其他都很一般般吧！【性价比】性价比就不说了直接满分  这么大的车裸车7w多块钱 去哪找？【为什么最终选择这款车？】其实购车前一直看中h6  但是资金有限（不想贷款）全身就10w  后来看了好多款  家里差点让买了宝骏560  和陆丰x7（家里支持资金）但是最后还是选择了s6 因为家里不喜欢比亚迪 这个名字（大家好多都懂的）说十几万宁愿买个CRV  不过我不喜欢日产（还是应人而异）【其他描述】|http://k.autohome.com.cn/spec/18563/view_1041472_1.html?st=184&piap=0 2088 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498388891|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 09:52:02|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=173&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498388918|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 09:52:02|2016年05月19日 发表了质量评价|2016年05月19日 发表了质量评价  质量   【行驶过程】  刹车时有异响-车辆前部  【内饰】  随车脚垫会滑动或污损       来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=155&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498388922|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 09:52:02|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=152&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498389051|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 09:52:02|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=61&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498389067|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 09:52:02|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=47&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498389100|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 09:52:02|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=24&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498406024|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-14 10:01:04|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=16&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498410001|Autohome_review|아반떼 AD(领动)|ZHO|2016-06-14 10:03:02|2016年06月02日 发表了口碑|来自：手机汽车之家  2016年06月02日 发表了口碑  口碑    《外观拉风 配置足够 整体性价比还是不错的。》           【最满意的一点】外观很拉风 现在路上还很少见 大轮毂。日间行车灯很高大上 自动头灯也很高端。中控台是软的 车内显示屏清晰度很高。倒车影像有随动辅助导线。很方便。车内音响很赞 我喜欢听音乐 完全满足我的要求。【最不满意的一点】后排不能放倒 这个真心很郁闷 这个放倒真的很难吗？这几天B柱内有异响 这还是新车呀 哎。。过几天去4s看看 希望不是啥大问题。另外胎噪确实大 我想跟轮胎大也有关系吧。悬挂还是有点硬 不过在接受范围内。【空间】空间同级别还是有优势的 中间无凸起。【动力】动力够用 现在用的eco模式【操控】转向精准 没啥虚位。【油耗】表显6 肯定是不准的 等下次油表亮再算算。【舒适性】还可以 家用够了。【外观】满意【内饰】做工还是比较好的 接缝均匀。【性价比】性价比高【为什么最终选择这款车？】同级别都看了 也试驾了 福克斯空间太小 科鲁兹都说油耗高 新英朗有点老气 卡罗拉没esp 思域根本没现车 看来看去家用也就韩系车了。【其他描述】换车的想法去年就有了 但是一直没有付诸行动 一是因为暂时有车开 二是今年上市新车多 想再等等 经常看论坛 心里已经有了几个备选 英朗 老表刚买的 开始觉得性价比很高 后来发现新旧差别很大 就pass了。福克斯外观不错 但是同事有好几辆 不想买一样的。k3性价比很高 优惠很大 但是新款感觉你没老款好看。看到最后就是领动了 配置高 外观拉风 总体性价比很高。|http://k.autohome.com.cn/spec/25701/view_1148059_1.html?st=43&piap=0 3959 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498416966|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-14 10:06:08|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=194&piap=0 657 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498480099|Autohome_review|뉴 보라(宝来)|ZHO|2016-06-14 10:42:01|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=220&piap=0 633 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498488313|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-14 10:47:13|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=197&piap=0 657 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498503149|365care|汽车|ZHO|2016-06-14 10:54:02|选一辆轿车很难吗？咱们看销量选肯定没错|选一辆轿车很难吗？咱们看销量选肯定没错_365关注网2016-06-14 09:43:00   来源：车早茶     点上方蓝字可加关注微信号：车早茶本文为车早茶原创文章 作者陈耀峰 转载请注明出处及作者2016年5月中国汽车销量已经出炉 经历了4月份的销量放缓之后 5月份的汽车整体销量趋向平稳 轿车市场方面 也还是平稳的态势。在榜单前十名中 合资品牌轿车依然一家独大 4月和5月榜单对比可见德系和美系车型销量持续火热。下面 茶哥就来给大家盘点一下5月份销量排名前十的轿车车型吧。>>>>第十名：科鲁兹5月份销量：16667辆茶哥辣评：在3月份排名15名的科鲁兹 此次挤掉起亚k3 杀入排行榜第十名 让人有点意外。不过科鲁兹也是款挺好的车 加上操控性好 外观也很耐看 排进前十也是有它的原因的。>>>>第九名：大众全新Polo5月份销量：16915辆茶哥辣评：诞生30年历经五代产品演变 总产量超过700万辆 并曾长期位居德国经济性小型车销量榜首 被称为德国大众的“神奇小子”。每次新款都吸引众多消费者选择 4月份排在轿车销量第14 这个月上升到第9。>>>>第八名：现代朗动5月份销量：18152辆茶哥辣评：朗动一直是8-10万区间的合资紧凑车的首选车型之一 纵使换代车型领动已经上市有一段时间 但它各方面都不算落后 再加上超高的性价比 领动想取代朗动估计还要很长时间。>>>>第七名：福特福睿斯4月份销量：21010辆茶哥辣评：福睿斯依然站稳在轿车销量的第七位 鸡蛋里面挑刺可能就要说比上月少卖1295辆 福睿斯源自福克斯平台 但定位比福克斯要低 它的热销证明了国人更在乎的是价格和空间 至于舒适度根本不是那么重要。>>>>第六名：大众速腾5月份销量：27988辆茶哥辣评：虽然跟上月比较 大众速腾下滑了一位 但速腾已经成为轿车销量榜前十的常客 直接原因肯定就是速腾的销量曲线没有走过山车 一直都较为稳定。可以看出它已经用实力在说服挑选它的消费者。>>>>第五名：日产轩逸5月份销量：28704辆茶哥辣评：说到轩逸 在日系车中算是销量的佼佼者 曾经也有人“埋怨”过轩逸变成街车 路上它的身影无处不在 这都要多得它的各方面都满足到国人 省油、舒适、空间大 而且毛病少 这样的车能不热销吗？>>>>第四名：丰田卡罗拉5月份销量：29318辆茶哥辣评：卡罗拉 身为全球销量第一的车型 但在国人心目中占比却不重 原因就应该不用多说了。但是推出了双擎版本后 卡罗拉的魅力就有所增加了。这也是今年长期能够活跃在销量榜前十内的一个原因。>>>>第三名：别克全新英朗5月份销量：30343辆茶哥辣评：这辆凯越平台的英朗 作为 “中国特供车”的表现非常出色 新款出来后 外形更好看 优惠更大 性价比更高 销量一直比较乐观。再加上凯越真正的换代车型威朗跟全新英朗的定位差距比较大 自然而然很多人都会选择买英朗。>>>>第二名：大众捷达5月份销量：30546辆茶哥辣评：当年老捷达积攒下来的优秀口碑 令到不少人为新捷达的情怀买单 所以销量表现也一直稳定 不过今年众多车型年轻化 捷达面临的竞争才刚刚开始。>>>>第一名：大众新朗逸5月份销量：36047辆茶哥辣评：朗逸在这个月比4月份销量多了1544辆 虽然离3月份的销量新高已经过了两个月 但他的销量还是坐稳在轿车销量排行榜的第一名 品牌魅力和实在的表现成为了它的吸睛点。茶哥总结：合资品牌再一个月占据了轿车销量排行榜的前十 虽然这两年自主品牌销量不断上升 但是如果要和传统的合资品牌更为正面的竞争估计还要加把劲 在各方面说服面临买车换车的消费者 要不然合资品牌在轿车领域的地位可能就更难挑战了。|http://www.365care.cn/2016/0614/3265146.html|2016-06-14
기타|2498505717|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 10:56:02|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=26&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498514401|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-14 11:02:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=193&piap=0 78 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498560793|Autohome_review|BYD S6(比亚迪S6)|ZHO|2016-06-14 11:27:12|2016年04月01日 发表了口碑|来自：汽车之家iPhone版  2016年04月01日 发表了口碑  口碑    《空间大就不用说了 没有之前担心的动力不足 感觉动力够用》           【最满意的一点】空间 配置 虽然2.0手豪（不想要天窗 应人而异）但是后期选装自装也是感觉很霸气 好多十多万的车都没有的配置  心里美滋滋～【最不满意的一点】目前就发现右后轮起步有点异响 但是说来也怪  每次到4s店就没有了 去了四五次都不响了 回家没几天又继续  好邪～【空间】前几天去了东北  （有贴） 后面气垫床谁俩人（178cm）没问题  还能装点东西～【动力】没有网上说的那么肉  我只想说只要舍得给油什么车都不肉【操控】开的还不错  就是刚开始开离合太高不习惯  现在习惯了 感觉很透  油门也挺灵活  （之前在部队开猛士） 开小六感觉 很棒【油耗】比预计要低可能跑长途的 以前市区差不多9个油还能接受 这次高速回来平均降到8.7 不管多少2.0这么大的车 只要不超十个油都能接受【舒适性】椅子倍舒服 以前猛士没法比  也不能比 不是一个级别 感觉比朋友的k3舒服多了！【外观】外观挺不错的  不过现在出来好的新车自然小六要逊色不少  不过自己折腾加装踏板 牛头杠 行李架 （准备换Q5大灯和仿宝马LED尾灯）【内饰】内饰除了座椅和方向盘很满意 其他都很一般般吧！【性价比】性价比就不说了直接满分  这么大的车裸车7w多块钱 去哪找？【为什么最终选择这款车？】其实购车前一直看中h6  但是资金有限（不想贷款）全身就10w  后来看了好多款  家里差点让买了宝骏560  和陆丰x7（家里支持资金）但是最后还是选择了s6 因为家里不喜欢比亚迪 这个名字（大家好多都懂的）说十几万宁愿买个CRV  不过我不喜欢日产（还是应人而异）【其他描述】|http://k.autohome.com.cn/spec/18563/view_1041472_1.html?st=185&piap=0 2088 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498571939|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-14 11:33:01|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=17&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498582692|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 11:39:01|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=177&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498582731|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 11:39:01|2016年05月19日 发表了质量评价|2016年05月19日 发表了质量评价  质量   【行驶过程】  刹车时有异响-车辆前部  【内饰】  随车脚垫会滑动或污损       来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=159&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498582737|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 11:39:01|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=156&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498582978|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 11:39:06|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=65&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498583030|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 11:39:06|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=51&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498583084|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 11:39:07|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=28&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498598292|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-14 11:47:32|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=198&piap=0 657 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498604603|sohu_auto|搜狐汽车 > 买车指导|ZHO|2016-06-14 11:50:01|选一辆轿车很难？看销量选肯定没错！|　　本文为车早茶原创文章 作者陈耀峰 转载请注明出处及作者 　　2016年5月中国汽车销量已经出炉 经历了4月份的销量放缓之后 5月份的汽车整体销量趋向平稳 轿车市场方面 也还是平稳的态势。在榜单前十名中 合资品牌轿车依然一家独大 4月和5月榜单对比可见德系和美系车型销量持续火热。下面 茶哥就来给大家盘点一下5月份销量排名前十的轿车车型吧。   　　>>>> 　　第十名：科鲁兹 　　5月份销量：16667辆  　　茶哥辣评：在3月份排名15名的科鲁兹 此次挤掉起亚k3 杀入排行榜第十名 让人有点意外。不过科鲁兹也是款挺好的车 加上操控性好 外观也很耐看 排进前十也是有它的原因的。 　　>>>> 　　第九名：大众全新Polo 　　5月份销量：16915辆  　　茶哥辣评：诞生30年历经五代产品演变 总产量超过700万辆 并曾长期位居德国经济性小型车销量榜首 被称为德国大众的“神奇小子”。每次新款都吸引众多消费者选择 4月份排在轿车销量第14 这个月上升到第9。 　　>>>> 　　第八名：现代朗动 　　5月份销量：18152辆  　　茶哥辣评：朗动一直是8-10万区间的合资紧凑车的首选车型之一 纵使换代车型领动已经上市有一段时间 但它各方面都不算落后 再加上超高的性价比 领动想取代朗动估计还要很长时间。 　　>>>> 　　第七名：福特福睿斯 　　4月份销量：21010辆 　　茶哥辣评：福睿斯依然站稳在轿车销量的第七位 鸡蛋里面挑刺可能就要说比上月少卖1295辆 福睿斯源自福克斯平台 但定位比福克斯要低 它的热销证明了国人更在乎的是价格和空间 至于舒适度根本不是那么重要。 　　>>>> 　　第六名：大众速腾 　　5月份销量：27988辆 　　茶哥辣评：虽然跟上月比较 大众速腾下滑了一位 但速腾已经成为轿车销量榜前十的常客 直接原因肯定就是速腾的销量曲线没有走过山车 一直都较为稳定。可以看出它已经用实力在说服挑选它的消费者。 　　>>>> 　　第五名：日产轩逸 　　5月份销量：28704辆  　　茶哥辣评：说到轩逸 在日系车中算是销量的佼佼者 曾经也有人“埋怨”过轩逸变成街车 路上它的身影无处不在 这都要多得它的各方面都满足到国人 省油、舒适、空间大 而且毛病少 这样的车能不热销吗？ 　　>>>> 　　第四名：丰田卡罗拉 　　5月份销量：29318辆  　　茶哥辣评：卡罗拉 身为全球销量第一的车型 但在国人心目中占比却不重 原因就应该不用多说了。但是推出了双擎版本后 卡罗拉的魅力就有所增加了。这也是今年长期能够活跃在销量榜前十内的一个原因。 　　>>>> 　　第三名：别克全新英朗 　　5月份销量：30343辆 　　茶哥辣评：这辆凯越平台的英朗 作为 “中国特供车”的表现非常出色 新款出来后 外形更好看 优惠更大 性价比更高 销量一直比较乐观。再加上凯越真正的换代车型威朗跟全新英朗的定位差距比较大 自然而然很多人都会选择买英朗。 　　>>>> 　　第二名：大众捷达 　　5月份销量：30546辆  　　茶哥辣评：当年老捷达积攒下来的优秀口碑 令到不少人为新捷达的情怀买单 所以销量表现也一直稳定 不过今年众多车型年轻化 捷达面临的竞争才刚刚开始。 　　>>>> 　　第一名：大众新朗逸 　　5月份销量：36047辆  　　茶哥辣评：朗逸在这个月比4月份销量多了1544辆 虽然离3月份的销量新高已经过了两个月 但他的销量还是坐稳在轿车销量排行榜的第一名 品牌魅力和实在的表现成为了它的吸睛点。 　　茶哥总结： 　　合资品牌再一个月占据了轿车销量排行榜的前十 虽然这两年自主品牌销量不断上升 但是如果要和传统的合资品牌更为正面的竞争估计还要加把劲 在各方面说服面临买车换车的消费者 要不然合资品牌在轿车领域的地位可能就更难挑战了。 　　买车用车不想被忽悠 　　关注微信号：车早茶   http://auto.sohu.com/********/n*********.shtml auto.sohu.com true 搜狐媒体平台  http://auto.sohu.com/********/n*********.shtml report 7419 本文为车早茶原创文章 作者陈耀峰 转载请注明出处及作者2016年5月中国汽车销量已经出炉 经历了4月份的销量放缓之后 5月份的汽车整体销量趋向平稳 轿车市场方面|http://auto.sohu.com/20160614/n454288927.shtml|2016-06-14
기타|2498648884|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-14 12:14:03|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=194&piap=0 78 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498651795|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-14 12:15:03|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=18&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498665814|Autohome_review|아반떼 AD(领动)|ZHO|2016-06-14 12:23:01|2016年06月02日 发表了口碑|来自：手机汽车之家  2016年06月02日 发表了口碑  口碑    《外观拉风 配置足够 整体性价比还是不错的。》           【最满意的一点】外观很拉风 现在路上还很少见 大轮毂。日间行车灯很高大上 自动头灯也很高端。中控台是软的 车内显示屏清晰度很高。倒车影像有随动辅助导线。很方便。车内音响很赞 我喜欢听音乐 完全满足我的要求。【最不满意的一点】后排不能放倒 这个真心很郁闷 这个放倒真的很难吗？这几天B柱内有异响 这还是新车呀 哎。。过几天去4s看看 希望不是啥大问题。另外胎噪确实大 我想跟轮胎大也有关系吧。悬挂还是有点硬 不过在接受范围内。【空间】空间同级别还是有优势的 中间无凸起。【动力】动力够用 现在用的eco模式【操控】转向精准 没啥虚位。【油耗】表显6 肯定是不准的 等下次油表亮再算算。【舒适性】还可以 家用够了。【外观】满意【内饰】做工还是比较好的 接缝均匀。【性价比】性价比高【为什么最终选择这款车？】同级别都看了 也试驾了 福克斯空间太小 科鲁兹都说油耗高 新英朗有点老气 卡罗拉没esp 思域根本没现车 看来看去家用也就韩系车了。【其他描述】换车的想法去年就有了 但是一直没有付诸行动 一是因为暂时有车开 二是今年上市新车多 想再等等 经常看论坛 心里已经有了几个备选 英朗 老表刚买的 开始觉得性价比很高 后来发现新旧差别很大 就pass了。福克斯外观不错 但是同事有好几辆 不想买一样的。k3性价比很高 优惠很大 但是新款感觉你没老款好看。看到最后就是领动了 配置高 外观拉风 总体性价比很高。|http://k.autohome.com.cn/spec/25701/view_1148059_1.html?st=42&piap=0 3959 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498707610|0797sf|汽车|ZHO|2016-06-14 12:47:17|选一辆轿车很难?看销量选肯定没错!|本文为车早茶原创文章 作者陈耀峰 转载请注明出处及作者2016年5月中国汽车销量已经出炉 经历了4月份的销量放缓之后 5月份的汽车整体销量趋向平稳 轿车市场方面 也还是平稳的态势。在榜单前十名中 合资品牌轿车依然一家独大 4月和5月榜单对比可见德系和美系车型销量持续火热。下面 茶哥就来给大家盘点一下5月份销量排名前十的轿车车型吧。>>>>第十名:科鲁兹5月份销量:16667辆茶哥辣评:在3月份排名15名的科鲁兹 此次挤掉起亚k3 杀入排行榜第十名 让人有点意外。不过科鲁兹也是款挺好的车 加上操控性好 外观也很耐看 排进前十也是有它的原因的。第九名:大众全新Polo5月份销量:16915辆茶哥辣评:诞生30年历经五代产品演变 总产量超过700万辆 并曾长期位居德国经济性小型车销量榜首 被称为德国大众的“神奇小子”。每次新款都吸引众多消费者选择 4月份排在轿车销量第14 这个月上升到第9。第八名:现代朗动5月份销量:18152辆茶哥辣评:朗动一直是8-10万区间的合资紧凑车的首选车型之一 纵使换代车型领动已经上市有一段时间 但它各方面都不算落后 再加上超高的性价比 领动想取代朗动估计还要很长时间。第七名:福特福睿斯4月份销量:21010辆茶哥辣评:福睿斯依然站稳在轿车销量的第七位 鸡蛋里面挑刺可能就要说比上月少卖1295辆 福睿斯源自福克斯平台 但定位比福克斯要低 它的热销证明了国人更在乎的是价格和空间 至于舒适度根本不是那么重要。第六名:大众速腾5月份销量:27988辆茶哥辣评:虽然跟上月比较 大众速腾下滑了一位 但速腾已经成为轿车销量榜前十的常客 直接原因肯定就是速腾的销量曲线没有走过山车 一直都较为稳定。可以看出它已经用实力在说服挑选它的消费者。第五名:日产轩逸5月份销量:28704辆茶哥辣评:说到轩逸 在日系车中算是销量的佼佼者 曾经也有人“埋怨”过轩逸变成街车 路上它的身影无处不在 这都要多得它的各方面都满足到国人 省油、舒适、空间大 而且毛病少 这样的车能不热销吗?第四名:丰田卡罗拉5月份销量:29318辆茶哥辣评:卡罗拉 身为全球销量第一的车型 但在国人心目中占比却不重 原因就应该不用多说了。但是推出了双擎版本后 卡罗拉的魅力就有所增加了。这也是今年长期能够活跃在销量榜前十内的一个原因。第三名:别克全新英朗5月份销量:30343辆茶哥辣评:这辆凯越平台的英朗 作为 “中国特供车”的表现非常出色 新款出来后 外形更好看 优惠更大 性价比更高 销量一直比较乐观。再加上凯越真正的换代车型威朗跟全新英朗的定位差距比较大 自然而然很多人都会选择买英朗。第二名:大众捷达5月份销量:30546辆茶哥辣评:当年老捷达积攒下来的优秀口碑 令到不少人为新捷达的情怀买单 所以销量表现也一直稳定 不过今年众多车型年轻化 捷达面临的竞争才刚刚开始。第一名:大众新朗逸5月份销量:36047辆茶哥辣评:朗逸在这个月比4月份销量多了1544辆 虽然离3月份的销量新高已经过了两个月 但他的销量还是坐稳在轿车销量排行榜的第一名 品牌魅力和实在的表现成为了它的吸睛点。茶哥总结:合资品牌再一个月占据了轿车销量排行榜的前十 虽然这两年自主品牌销量不断上升 但是如果要和传统的合资品牌更为正面的竞争估计还要加把劲 在各方面说服面临买车换车的消费者 要不然合资品牌在轿车领域的地位可能就更难挑战了。     网友评论|http://www.0797sf.com/2016-06-14/3267028.html|2016-06-14
기타|2498721539|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-14 12:57:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=199&piap=0 657 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498750812|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-14 13:15:04|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=195&piap=0 78 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498785199|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-14 13:36:01|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=201&piap=0 657 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498815106|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-14 13:54:03|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=19&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498826110|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 14:01:02|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=179&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498826155|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 14:01:02|2016年05月19日 发表了质量评价|2016年05月19日 发表了质量评价  质量   【行驶过程】  刹车时有异响-车辆前部  【内饰】  随车脚垫会滑动或污损       来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=161&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498826162|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 14:01:02|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=158&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498826420|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 14:01:02|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=67&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498826466|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 14:01:02|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=53&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498826542|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 14:01:02|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=29&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498850937|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-14 14:16:01|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=204&piap=0 657 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498851171|Autohome_review|뉴 보라(宝来)|ZHO|2016-06-14 14:16:01|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=222&piap=0 633 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498853032|Autohome_review|BYD S6(比亚迪S6)|ZHO|2016-06-14 14:17:01|2016年04月01日 发表了口碑|来自：汽车之家iPhone版  2016年04月01日 发表了口碑  口碑    《空间大就不用说了 没有之前担心的动力不足 感觉动力够用》           【最满意的一点】空间 配置 虽然2.0手豪（不想要天窗 应人而异）但是后期选装自装也是感觉很霸气 好多十多万的车都没有的配置  心里美滋滋～【最不满意的一点】目前就发现右后轮起步有点异响 但是说来也怪  每次到4s店就没有了 去了四五次都不响了 回家没几天又继续  好邪～【空间】前几天去了东北  （有贴） 后面气垫床谁俩人（178cm）没问题  还能装点东西～【动力】没有网上说的那么肉  我只想说只要舍得给油什么车都不肉【操控】开的还不错  就是刚开始开离合太高不习惯  现在习惯了 感觉很透  油门也挺灵活  （之前在部队开猛士） 开小六感觉 很棒【油耗】比预计要低可能跑长途的 以前市区差不多9个油还能接受 这次高速回来平均降到8.7 不管多少2.0这么大的车 只要不超十个油都能接受【舒适性】椅子倍舒服 以前猛士没法比  也不能比 不是一个级别 感觉比朋友的k3舒服多了！【外观】外观挺不错的  不过现在出来好的新车自然小六要逊色不少  不过自己折腾加装踏板 牛头杠 行李架 （准备换Q5大灯和仿宝马LED尾灯）【内饰】内饰除了座椅和方向盘很满意 其他都很一般般吧！【性价比】性价比就不说了直接满分  这么大的车裸车7w多块钱 去哪找？【为什么最终选择这款车？】其实购车前一直看中h6  但是资金有限（不想贷款）全身就10w  后来看了好多款  家里差点让买了宝骏560  和陆丰x7（家里支持资金）但是最后还是选择了s6 因为家里不喜欢比亚迪 这个名字（大家好多都懂的）说十几万宁愿买个CRV  不过我不喜欢日产（还是应人而异）【其他描述】|http://k.autohome.com.cn/spec/18563/view_1041472_1.html?st=187&piap=0 2088 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498854847|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-14 14:18:02|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=21&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498921085|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-14 14:56:01|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=205&piap=0 657 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2498985287|Autohome_review|뉴 보라(宝来)|ZHO|2016-06-14 15:30:02|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=223&piap=0 633 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499040586|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-14 16:01:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=206&piap=0 657 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499041502|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-14 16:01:07|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=23&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499060506|Autohome_review|뉴 보라(宝来)|ZHO|2016-06-14 16:11:02|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=224&piap=0 633 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499107488|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-14 16:36:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=207&piap=0 657 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499110892|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-14 16:38:02|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=24&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499173945|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-14 17:10:04|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=26&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-14
其他媒体|2499188996|difang CN|地方频道 > 滚动读报|ZHO|2016-06-14 17:17:02|2016ctcc转战珠海 新k3势头不减再获冠军|6月5日 2016年ctcc中国房车锦标赛移师广东珠海。在首站取得惊艳成绩的东风悦达起亚势头不减 借助实力强劲的新k3再下一城 拿下珠海站超级杯1.6t组厂商杯冠军。在目前已经结束的两站赛事中 叶弘历、詹家图、张志强、林立峰所组成的王牌车队之所以能所向披靡包揽超级杯1.6t组厂商杯冠军 新k3的作用功不可没。新k3在5月也取得近1.5万台的骄人业绩 位列细分市场领先位置 可谓名利双收。据悉 ctcc的战火接下来将席卷上海、韩国全罗道等城市 相信新k3也会愈战愈勇 带来更加精彩的表现 让我们拭目以待。（起亚）|http://difang.gmw.cn/newspaper/2016-06/14/content_113217573.htm|2016-06-14
기타|2499194724|SINA_auto|导购 > 车型导购|ZHO|2016-06-14 17:20:01|几款值得买的8-10万元家用SUV！|　　近几天有不少朋友留言问小编“8—10万的SUV有哪些值得买？”首先小编在这里先感谢一下各位看观们对《汽车大观》的支持 小编的膝盖已经献上。好了 咱们说正事 小编看到留言那以后就开始苦（百）苦（度）思（一）索（下） 目前市场上有哪些8—10万范围内的SUV 经过小编的一番搜索 在这里小编就为各位看观们推荐几款值得买的8—10万元的家用SUV。　　帝豪GS　　售价7.78-10.88万元　　5月4日 吉利汽车宣布吉利帝豪GS上市 新车共推出1.3T和1.8L两种排量总计11款车型 官方指导价为7.78万-10.88万元。　　帝豪GS在延续吉利全新家族式设计语言的基础上 融入了更多当下年轻人喜爱的现代时尚元素 动感前卫的跨界造型、精致时尚的内饰、越级安全配置等 都彰显了帝豪GS年轻时尚的跨界风格与精致品质。　　车身的长宽高分别为4440/1833/1560mm 轴距达到2700mm。ACC自适应巡航系统、预碰撞安全系统、ESP车身电子稳定系统、TPMS智能胎压监测系统、电子驻车EPB+AUTOHOLD、GSG智能启停系统以及EPS电动随速助力转向在内的丰富的配置加上7.78-10.88万元的售价 使得该车具有相当高的性价比。　　总结：　　优点： 　　1、漂亮的外观以及超控台做工精良　　2、不错的动力　　3、良好的操控和隔音效果　　4、低油耗　　5、良好的舒适性　　缺点：  　　1、后备箱空间略小　　2、天窗无法打开　　3、后梁非独立　　推荐指数：★★★★☆（四星半）　　长安CS75　　qichedaguan　　售价9.28—15.28万元　　3月22日 2016款长安CS75全新升级上市 官方指导价仅9.28万元起。2016款CS75新增的车头灵动双环形LED日行灯 以及车尾炫彩点亮式尾灯。全系车型由原来2014款的杆式天线升级为鲨鱼鳍天线 并新增双边排气布局。CS75的轴距达到2700mm 使得车辆拥有超大的空间尺度。　　CS75的安全配置有ESP系统 全车6安全气囊、ESC、AUTO-HOLD电子驻车系统、BLIS并线辅助系统、盲区监测系统、胎压监测系统、EPB电子驻车系统等。　　在动力上 2016款CS75搭载D20VVT发动机 最大功率116KW 最大扭矩200N.m 匹配高效 6速手动变速器。　　舒适性上 2016款长安CS75的长/宽/高仍旧保持4650mm/1850mm/1705mm 轴距为2700mm 具有大尺寸的肩部空间、肘部空间和臀部空间。　　长安CS75的配置相当丰富 包括NVH超静音、EPS电动助力精准操控、全自动空调配置、皮质电动6向可调节座椅+加热功能、智能无钥匙启动、搭载全面升级版 in Call智能车载互联系统、EPB电子手刹、无钥匙进入、一键启动、一键升降、后排空调出风口等功能。　　总结：　　优点：　　1、静音效果好　　2、外观时尚大气、空间大　　3、动力够用　　4、舒适度较高　　5、配置齐全、性价比高　　缺点：　　1、悬挂偏硬　　2、油耗高　　3、风噪较大　　4、座椅相对较硬　　推荐指数：★★★★☆（四星半）　　宝骏560　　qichedaguan　　售价7.68-9.08万元　　作为宝骏推出的首款紧凑型SUV车型 这款车主销车型价格在8万元左右 相对其它自主品牌SUV拥有强大竞争力。就产品本身来说 空间非常宽大 外观内饰设计颇为时尚精致。　　宝骏560在外观方面采用了宝骏家族式的盾形前进气格栅 略微修饰的镀铬装饰进气格栅并不显眼但足够提气。在灯光的使用上 宝骏560采用了LED日行灯和转向灯 并为大灯使用了透镜 整体上颇具动感。同时尾灯同样使用了LED光源 在功能方面 倒车雷达为全系标配 中高配还配有倒车影像。　　宝骏560轴距2750mm的  1.8L自然吸气发动机 最大功率101kW 峰值扭矩186N/m。动力不弱 也够给劲儿。配置上面也比较丰富 560带有用户记忆模式的8英寸触摸式大屏 集GPS、蓝牙、广播、CD、手机映射等功能于一身 车子还配置了一键启动、多功能方向盘、定速巡航等等都很实用。　　总结：　　优点： 　　1、空间大、坐姿高　　2、操控性 风噪、胎噪比较好　　3、油耗低　　4、底盘较稳　　缺点： 　　1、动力不足 提速慢　　2、灯光较弱　　3、导航不太准、收音机效果差、外循环空调制冷效果差　　推荐指数：★★★☆（三星半）　　大迈X5　　qichedaguan　　售价7.39-10.89万元　　大迈X5配置丰富 乘坐和储物空间也能很好满足一般家庭需求 大迈X5的外观很有质感。　　众泰大迈X5长宽高依次为4527/1836/1682mm 轴距达到了2680mm 最小离地间隙为180mm 各项数据在国内同级车型中都综合领先 对于家用来说空间绝对够用。　　T型布局的中控台少了很多复杂的设计与配饰 黑色的主题颜色让人感觉十分干练。内饰同样采用了大量的平直硬朗的线条 配合钢琴烤漆和亮条元素 极具时尚感。　　在安全性配置部分 新车全系标配防眩目内后视镜、ISOFIX儿童安全座椅固定接口、前排双安全气囊、主驾驶安全带未系提醒、电子手刹、ABS+EBD、后倒车雷达等。　　顶配车型则会增配前排侧安全气囊、头部气帘、ESC等。在外观和内饰配置方面 大迈X5将会全系标配LED日间行车灯、后雾灯、LED尾灯、电动调节外后视镜等。　　在舒适及科技配置部分 大迈X5会标配真皮多功能方向盘、四门电动车窗、遥控停车、遥控中央门锁等。高配车型则还会配备全景天窗、一键启动/无钥匙进入、8英寸液晶显示屏、倒车影像等。顶配车型则还会配备自动恒温空调。　　大迈X5车型搭载三菱1.5T涡轮增压发动机 并配备5挡手动变速器。三菱1.5T涡轮增压发动机采用MIVEC进气连续可变气门正时机构 全铝材质使整个发动机更加轻量化 加上性能优良的增压器 最大功率达到110kW/6000rpm 最大扭矩195Nm/****-****rpm 可以为大迈X5提供动力。与之匹配5速手动和CVT无极变速箱。　　8万最低配版本就能够开回家 驾驶轻松 配置丰富 够用的动力 这几个有点使得大迈X5是一款不错的家用车。　　总结：　　优点：　　1、外观大气、内饰用料考究　　2、滤震舒适、空间大　　3、配置丰富、性价比高　　4、油耗低　　缺点： 　　1、非顶配车型全景天窗不能打开　　2、隔音效果一般　　3、涡轮介入前动力较差　　4、方向盘只有两项调节　　5、变速箱顿挫比较明显　　推荐指数：★★★☆（三星半）　　瑞虎5 　　qichedaguan　　售价8.99-15.09万元　　瑞虎5有着时尚大气的外观 经济省油的动力 是一款具有高适应性的家庭SUV。瑞虎5的安全性 多功能性和舒适性是它最大的亮点。　　安全性： 车身关键部位采用了屈服强度在1000MPa以上的高强度钢材。而且从中配的车开始导航就有定速巡航 超速报警。 顶配的车身更含有博士9.0的ESP7位一体的车身安全系统：ABS、EBD、TCS、DTC、HHC、ESM、HBA。　　多功能性 就是指车身的各种路面通过性 它的底盘满载里地间隙是168mm 轮胎规格是225。　　总结：　　优点：　　1、操控灵活简便 整体舒适　　2、底盘高　　3、时尚大气的外观时尚大气　　4、配置丰富 性价比高　　缺点：　　1、后备箱空间较小　　2、天窗偏小　　3、动力不足　　4、噪音较大　　推荐指数：★★★★（四星）　　（来源：汽车大观）|http://auto.sina.com.cn/mp/g/2016-06-14/detail-ifxszfak3740424.shtml|2016-06-14
기타|2499207068|Autohome_review|아반떼 AD(领动)|ZHO|2016-06-14 17:27:31|2016年06月02日 发表了口碑|来自：手机汽车之家  2016年06月02日 发表了口碑  口碑    《外观拉风 配置足够 整体性价比还是不错的。》           【最满意的一点】外观很拉风 现在路上还很少见 大轮毂。日间行车灯很高大上 自动头灯也很高端。中控台是软的 车内显示屏清晰度很高。倒车影像有随动辅助导线。很方便。车内音响很赞 我喜欢听音乐 完全满足我的要求。【最不满意的一点】后排不能放倒 这个真心很郁闷 这个放倒真的很难吗？这几天B柱内有异响 这还是新车呀 哎。。过几天去4s看看 希望不是啥大问题。另外胎噪确实大 我想跟轮胎大也有关系吧。悬挂还是有点硬 不过在接受范围内。【空间】空间同级别还是有优势的 中间无凸起。【动力】动力够用 现在用的eco模式【操控】转向精准 没啥虚位。【油耗】表显6 肯定是不准的 等下次油表亮再算算。【舒适性】还可以 家用够了。【外观】满意【内饰】做工还是比较好的 接缝均匀。【性价比】性价比高【为什么最终选择这款车？】同级别都看了 也试驾了 福克斯空间太小 科鲁兹都说油耗高 新英朗有点老气 卡罗拉没esp 思域根本没现车 看来看去家用也就韩系车了。【其他描述】换车的想法去年就有了 但是一直没有付诸行动 一是因为暂时有车开 二是今年上市新车多 想再等等 经常看论坛 心里已经有了几个备选 英朗 老表刚买的 开始觉得性价比很高 后来发现新旧差别很大 就pass了。福克斯外观不错 但是同事有好几辆 不想买一样的。k3性价比很高 优惠很大 但是新款感觉你没老款好看。看到最后就是领动了 配置高 外观拉风 总体性价比很高。|http://k.autohome.com.cn/spec/25701/view_1148059_1.html?st=45&piap=0 3959 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499229320|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 17:38:05|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=182&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499229367|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 17:38:05|2016年05月19日 发表了质量评价|2016年05月19日 发表了质量评价  质量   【行驶过程】  刹车时有异响-车辆前部  【内饰】  随车脚垫会滑动或污损       来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=164&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499229370|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 17:38:05|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=161&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499229511|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 17:38:05|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=70&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499229531|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 17:38:05|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=56&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499229561|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 17:38:05|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=33&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499235320|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-14 17:41:04|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=210&piap=0 657 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499266022|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-14 17:56:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=199&piap=0 78 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499287063|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-14 18:07:52|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=27&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499381413|SINA_auto|导购 > 车型导购|ZHO|2016-06-14 18:57:02|16万起 高性价比大空间中型车这些划算|　　现如今 车型越来越多 自然竞争就越来越激烈 无论是在哪个级别。就中级车而言 很多合资车型的价格都已经下探到20万以下了 这也让很多预算在20以内的消费者有了更多的一个选择 所以今天就给大家介绍几款20以下就可以落地的中级车。　　上汽通用雪佛兰-迈锐宝　　指导价：16.49-19.99万元　　推荐车型：1.6T 自动豪华版秒车价 配置  图库  视频  口碑  经销商迈锐宝 16.49万-19.99万元询价　　迈锐宝多年积累起来的用户口碑还是很不错的 改款后的外观和内饰也更能取悦到国内年轻消费者。内饰在舒适度上得到一定提高 比同级别采用了更高级一些的皮革面料。但是空间仍然是个软肋 虽然算不上局促 但是相比起其他的中级车而言 后排空间仍有可提升的空间。　　在推荐车型上的配置算比较丰富 刹车辅助 车身稳定控制 倒车影像 自动大灯等很实用的配置基本配备。并且由于是1.6T车型所以可以享购置税减半政策 性价比还是不错的。　　广汽本田-雅阁　　指导价：16.98-23.78万　　推荐车型：2.0L 豪华版　　雅阁以往给人的感觉都一种比较老气稳重的感觉 但改款之后雅阁里里外外都“翻新”了一遍 除了外观更加年轻时尚之外 配置上也增加了不少 基本是做到了加量不加价的地步了。　　除了加入了苹果CarPlay和Honda SENSING智能辅助系统等科技配置之外 上坡辅助 自动驻车 倒车影像等日常比较常用到的都有配备。虽然取代V6的2.0L和2.4L发动机没有V6那么大魅力 但是油耗还是有所降低。　　东风悦达起亚-K5　　指导价：15.98-23.98万　　推荐车型：1.6T 自动LUXURY　　起来K5还是保持着它那一贯的设计风格 说他运动吧 好像不对 说他商务也好像不太对 也许这就是所谓的“韩国欧巴”。内饰的面板质地和做工上有着比较明显的进步 触感比较舒服。　　起亚K5的配置也还算是丰富 除了只有顶配车型才有的自动驻车 胎压监测 全景天窗等一些配置之外 其他车型都有配备车身稳定控制 刹车辅助等一些安全实用的配置。新增的1.6T发动机替代了原来的2.4L发动机 搭配双离合 动力输出平顺 提速也够快。同样1.6T车型可享购置税减半。　　总结：三款车都来自不同的派系 各自有着各自特点 迈锐宝有品质和口碑 雅阁价格更加亲民且不减“料” K5相对均匀一些 可以说三款车的群体不尽相同 而你是属于哪一个呢？|http://auto.sina.com.cn/mp/g/2016-06-14/detail-ifxszfak3785688.shtml|2016-06-14
기타|2499431480|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-14 19:25:03|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=28&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499460885|SINA_auto|新车 > 谍照|ZHO|2016-06-14 19:44:01|一汽大众新捷达外观升级|　　今年年初一汽-大众公布了2016年“发轫”计划 除大众品牌年销量将冲击130万辆目标之外 在产品方面还将推出多款新车型 根据大众汽车此前的规划 未来将投产排量为1.5升的发动机 并在旗下车型使用。我们获得了一组新款捷达车型谍照 新车外观方面较现款车型进行细节调整 同时将有望搭载最新的1.5升自然吸气发动机 燃油经济性表现突出。　　新款捷达在外观整体方面与现款车型基本相同 仅有几处细节进行微调。根据谍照来看 新车局部位置进行了伪装 因此有望在大灯组及前格栅上增加全新设计的装饰条 车身侧面增加防擦条 同时后杠也有望做出修改 尾灯则采用LED光源 效果较现款车型提升明显。　　现款捷达搭载1.4升、1.4T和1.6升三款发动机 其中1.4升发动机最大输出功率为66千瓦 1.4T发动机最大输出功率为96千瓦 1.6升发动机最大输出功率为81千瓦；三款发动机百公里油耗分别为5.9升、5.8升和6升。与现搭载的三款发动机相比 新增的1.5升发动机比1.4升发动机动力更好 和1.6升发动机动力持平 略逊于1.4T发动机。但燃油经济性上 1.5升发动机百公里油耗为5.7升 比上述三款发动机表现更为出色。　　动力方面与同级别车型相比 科鲁兹搭载的1.5升自然吸气发动机最大输出功率为84千瓦 峰值扭矩为146牛米 综合百公里油耗为6.2升。两车相比后 可以看到新款捷达1.5升发动机动力表现虽略逊于科鲁兹 但燃油经济性新款捷达比科鲁兹低0.5升。整体来看 拥有售价、燃油经济性等优势的新款捷达市场竞争力将进一步提升。　　现款捷达搭载1.6升发动机的车型 在价格当中包括了5%的消费税以及17%的增值税 在换装了更小排量的1.5升发动机之后对应税率为3% 下调了2个百分点 以目前8.5万元左右的售价计算 消费税若下降2个百分点相当于1700元左右。   视频加载中 请稍候...     自动播放            play 捷达宝来质惠版超值上市    向前 向后|http://auto.sina.com.cn/newcar/d/2016-06-14/detail-ifxszfak3806298.shtml|2016-06-14
기타|2499478437|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-14 19:54:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=200&piap=0 78 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499485837|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-14 19:58:03|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=30&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499509862|Autohome_review|아반떼 AD(领动)|ZHO|2016-06-14 20:13:01|2016年06月02日 发表了口碑|来自：手机汽车之家  2016年06月02日 发表了口碑  口碑    《外观拉风 配置足够 整体性价比还是不错的。》           【最满意的一点】外观很拉风 现在路上还很少见 大轮毂。日间行车灯很高大上 自动头灯也很高端。中控台是软的 车内显示屏清晰度很高。倒车影像有随动辅助导线。很方便。车内音响很赞 我喜欢听音乐 完全满足我的要求。【最不满意的一点】后排不能放倒 这个真心很郁闷 这个放倒真的很难吗？这几天B柱内有异响 这还是新车呀 哎。。过几天去4s看看 希望不是啥大问题。另外胎噪确实大 我想跟轮胎大也有关系吧。悬挂还是有点硬 不过在接受范围内。【空间】空间同级别还是有优势的 中间无凸起。【动力】动力够用 现在用的eco模式【操控】转向精准 没啥虚位。【油耗】表显6 肯定是不准的 等下次油表亮再算算。【舒适性】还可以 家用够了。【外观】满意【内饰】做工还是比较好的 接缝均匀。【性价比】性价比高【为什么最终选择这款车？】同级别都看了 也试驾了 福克斯空间太小 科鲁兹都说油耗高 新英朗有点老气 卡罗拉没esp 思域根本没现车 看来看去家用也就韩系车了。【其他描述】换车的想法去年就有了 但是一直没有付诸行动 一是因为暂时有车开 二是今年上市新车多 想再等等 经常看论坛 心里已经有了几个备选 英朗 老表刚买的 开始觉得性价比很高 后来发现新旧差别很大 就pass了。福克斯外观不错 但是同事有好几辆 不想买一样的。k3性价比很高 优惠很大 但是新款感觉你没老款好看。看到最后就是领动了 配置高 外观拉风 总体性价比很高。|http://k.autohome.com.cn/spec/25701/view_1148059_1.html?st=44&piap=0 3959 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499537727|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-14 20:29:03|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=201&piap=0 78 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499561055|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 20:43:01|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=185&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499561133|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 20:43:01|2016年05月19日 发表了质量评价|2016年05月19日 发表了质量评价  质量   【行驶过程】  刹车时有异响-车辆前部  【内饰】  随车脚垫会滑动或污损       来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=167&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499561147|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 20:43:01|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=164&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499561547|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 20:43:02|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=73&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499561583|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 20:43:02|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=59&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499561643|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 20:43:02|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=36&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499563046|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-06-14 20:44:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=208&piap=0 657 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499588059|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-14 20:59:03|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=202&piap=0 78 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499695775|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-14 22:03:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=203&piap=0 78 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499720585|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-14 22:17:01|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=29&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499743075|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 22:30:01|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=74&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499743099|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 22:30:01|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=60&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499743152|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 22:30:01|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=38&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499815014|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-14 23:16:44|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=204&piap=0 78 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499850262|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 23:38:01|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=75&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499850315|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 23:38:01|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=61&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499850387|Autohome_review|K3(起亚K3)|ZHO|2016-06-14 23:38:01|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=39&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-14
기타|2499874169|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-14 23:53:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=205&piap=0 78 0 0 2 0 0 0 0 0 1|2016-06-14
其他社区|1594767257|360doc|最新文章|ZHO|2015-01-04 17:53:02|30年代国军制式武器的优化配置方案（最新修改版）|30年代国军制式武器的优化配置方案（最新修改版）（总论）20世纪30年代 日本侵略中国的脚步日益临近。国民政府在德国顾问的帮助指导下 开始了整军计划 核心就是建立兵工装备体系和统一军队编制。在抗战爆发前 整军取得了一定的成效 并对抗战初期的战局发挥了积极作用。但是 无论是国民政府的军队领导人还是德国顾问 都存在时代的局限 对制式武器的选择存在一定不足 影响了作战效果。本文讨论的内容就是为抗战时期的中国军队选择最为合适的陆军制式武器 从而能在抗日战场上发挥出最大的战斗力。这种假想绝不是凭空胡编乱造 给国军装备一大堆先进武器 那样就太没有意义了。本文所有的论述都建立在20世纪30年代前期和中期的时代背景 仿制武器都是中国当时的工业水平所能生产的 进口武器都是当时国外已经存在并且适合中国国情的 绝对不会出现超越时代的先进武器 也不会突破当时中国的所能够达到的生产能力（或许稍微提高一点）。当然 我们现在讨论这些事 是基于几十年来的经验总结 掌握了前人所不能获取的大量信息。因此 我并无苛求前人做得不好的意思 只是想探讨和真实的历史相比 能否有更为科学的陆军制式武器规划 会达到怎么样的效果 以为后人借鉴。欢迎各位网友一同讨论指正 不过有几点要提请各位网友注意。1. 关于本文的主题：本文是一个技术贴 主要讨论装备方面的问题。我也知道30年代的国府和国军存在太多的问题 指挥系统 人员训练 动员能力 后勤保障等等 不客气地说 我比这里大多数人认识得要深刻许多。不过这些问题需要另外专门撰文论述 不可能在一篇文章内面面俱到。所以请网友们在发言前注意 不要离题太远了。2. 关于年代背景：本文说的很清楚 年代背景是30年代初期和中期 更准确地说是1936年之前。所以二次大战中才出现的武器 比如英国斯登冲锋枪 苏俄14.5mm反坦克枪 美国巴祖卡火箭筒之类的武器 各位网友就不要讨论了。请切记这一点。3. 关于国军制式武器的装备范围：当时中国还没有形成统一 工业能力也无法支持全面换装 这是客观事实。我从来没指望能在短期内实现全面换装 这些设想中的制式武器 最多也就装备少量中央军的精锐部队 其他部队还是要长时间使用各种老式杂牌武器。但对于国府来说 至少要给兵工体系设定一个基准目标 逐步调整 朝这个方向去努力。然后在战争过程中 杂牌武器慢慢损耗 新出厂的武器都是一个规格 逐渐地 制式统一就形成了。有一个标准 总比没有标准 仍然五花八门各自为政好吧？而且我提出的这个标准不是高不可攀 是可以实现的 装备少量精锐部队财政上也负担得起。4. 关于备选方案：   有些轻武器装备可以有不同的选择 也是很不错的配置。因此 我还设计了一套备用方案。备选方案的配置从战术性能上来说不是最优 但却是对工业能力要求相对较低 对30年代现存装备改动最小 比较省事的。可以供网友参考比较。5. 关于仿制和进口的区分：基于30年代民国的工业能力 想实现所有制式武器全部国产化是绝对不可能的 有限的工业资源和技术只能保证一些最基本的步兵武器。所以一些装备还只能靠少量进口。这就需要区分哪些可以仿制 哪些需要进口。我的观点是步枪、轻重机枪、手枪、冲锋枪、迫击炮和山炮是应该自产的；野炮、榴弹炮、高射炮、反坦克炮和大口径机枪就只能进口。请网友在讨论时先看清楚仿制和进口的设定 不要先下结论说某某武器造不出来。可能这某某武器本来就是应该进口的。（一）步枪弹步枪弹是所有弹药中影响面最广的一种 涉及到每个一线步兵。步枪弹的选择直接关系到步兵战斗力的发挥 也决定了步枪和机枪的制式 必须慎重考虑。（1）30年代各种步枪弹的优缺点分析20世纪初到抗战爆发为止 中国军事领域受德国和日本的影响很大 因此国内使用的步枪弹主要也是以德式和日式为主 德国7.92×57mm毛瑟步枪弹最多 日本6.5×50mm有坂步枪弹其次。其他很多种类的枪弹 如苏联7.62mm 莫辛-纳甘枪弹、奥地利8mm曼利夏步枪弹、意大利6.5mm卡尔卡诺步枪弹、英国0.303英寸李恩菲尔德步枪弹、法国8mm勒伯尔步枪弹等 国内都有使用 但装备数量都比较少。直到抗战后期 随着美国援助物资的到达 斯普林菲尔德0.30-06步枪弹的使用有所增加 但仍然不及德、日两种子弹普遍。近年来 随着网络普及 特别是军事玄幻小说兴起 各种以讹传讹的说法流传开来 给人们造成不少错觉。仿佛7.92×57mm毛瑟步枪弹和中正式步枪的组合 完全克制了6.5×50mm有坂步枪弹和三八式步枪的组合 抗战时中国军队的轻武器优于日本军队。实际上 7.92mm毛瑟步枪弹并非完美无缺 6.5mm有坂步枪弹也不是人们想像的那么差。7.92mm毛瑟步枪弹的优点是威力大 杀伤效果好 缺点是全弹的尺寸和质量都比较大 后坐力太大。基本上 当时流行的全威力枪弹 如7.92mm毛瑟步枪弹、斯普林菲尔德0.30-06步枪弹和苏联7.62mm 莫辛-纳甘枪弹都有类似的特点。口径在7.5～8mm之间 枪口功能在3500J~4000J之间。这类枪弹的远距离存能好 更适合作为机枪子弹 用于远距离火力压制；而作为步枪子弹 则显得威力过剩。7.92mm毛瑟步枪弹的后坐力对于身长体壮的欧美人种还能承受 对于个头普遍矮小一些的东亚人种而言就显得太大了。当时中国士兵普遍营养不良 身体瘦弱 尤其是对新兵而言 一下子使用这种全威力枪弹 很难控制好枪支。再加上当时中国军工生产能力薄弱 军队实弹训练少 没有机会去慢慢适应强大的后坐力。最终造成的后果就是士兵在战斗中控制不好步枪 射击精度不佳 子弹的杀伤力再大 打不准又有什么用？同时 在大规模战争时期 参战部队往往要持续作战好几天得不到休息 过大的后坐力很容易导致士兵疲劳 体力迅速下降 从而影响部队的持续作战能力。6.5mm有坂步枪弹的优点是射击精度高 后坐力小 缺点是远距离停止作用偏小。经过网络的渲染 人们对该弹的印象就是杀伤力小 容易形成贯通伤 毫无可取之处。其实这种理解并不全面 有坂弹容易穿透人体 并不是子弹本身的问题 而是发射该弹的三八式步枪枪管膛线缠距过短 子弹出膛转速过高引起的。所谓“一枪两个眼”的情况也不是很常见 只是概率高一些而已 不能把特例误认为普遍现象。后期经过改进 有坂弹的杀伤力明显有提高 太平洋战场上的美军调查报告中对该弹的评价就很好。有坂步枪弹后坐力小 有利于提高射击水准 特别对训练新兵很有帮助 减少其恐惧感 能很快掌握步枪使用要领。针对当时中国士兵缺乏训练的情况 实在是很有意义的。当时世界上采用6.5mm口径子弹的国家也不少 比如意大利使用的6.5×52mm卡尔卡诺步枪弹、荷兰／罗马尼亚使用的6.5×54mmR曼利夏步枪弹、瑞典使用的6.5×55mm毛瑟步枪弹等 其中以瑞典6.5mm毛瑟步枪弹性能最佳。这些6.5mm口径的枪弹枪口动能都在2500J～3000J之间 如果用于机枪火力压制 的确存在远距离停止作用偏小的缺点。但在用于步枪时 只要其威力能够满足在一定距离上精确射杀目标的要求 就已经足够了。后来发展的7.92×33mm和7.62×39mm等中间威力步枪弹的枪口动能都只有2000J上下 却很少听到有人说它们不行 因为它们的威力已经够用了。（2）采用7×57mm步枪弹适合中国战场的需要总的来说 枪口动能在3500J以上不适合做步枪弹 3000J以下不适合做机枪弹。如果要实现步机枪弹统一 就需要有一种性能平衡的子弹 既有较小的后坐力 又有较大的杀伤力 枪口动能在3000J～3500J之间。考虑到当时中国的工业水平 不可能设计全新的弹药 只能在当时已有的子弹中选择一种最符合上述要求的型号仿制 7×57mm毛瑟步枪弹无疑是最优选择。该型子弹由于最早为西班牙军队所装备 俗称西班牙毛瑟弹 实际上德国、比利时、捷克等都生产过 以比利时产量最大。拉美国家使用比较广泛 包括哥伦比亚、巴西、委内瑞拉、智利、墨西哥、多米尼加等。网上搜索到的关于该弹的数据多半是早期的圆头弹 事实上该弹在1913年已改为尖头弹。《金属与火焰的回忆：二战军用枪弹全接触》一文中就有图片。7×57mm毛瑟步枪弹的枪口功能约为3300J 弹头设计合理 初速高 后坐力较小 杀伤力较大 精度也很好 平衡兼顾了步枪和机枪两种需求。而且它的弹壳与的7.92×57mm步枪弹的弹壳基本相同 只是弹头收口处更小些。鉴于国内各兵工厂生产7.92×57mm步枪弹的经验较多 工艺设备调整量也不大 因此很容易大量生产。从性能和生产能力这两方面结合来看 7×57mm毛瑟步枪弹都很适合抗战时期中国军队的需求。（3）圆头弹和尖头弹的差异一定会有网友提出 从清末开始 中国的弹药种类已经很多 其中的主流枪弹又一直是德国7.92mm毛瑟步枪弹 改用一种新口径的弹药会增加兵工生产和后勤补给的困难 还是用7.92mm毛瑟步枪弹为佳。这种看法其实忽略了一个关键点 清末到30年代之前 中国各大兵工厂造的7.92mm毛瑟步枪弹几乎都是圆头弹 而不是尖头弹！圆头弹已经落后于时代 新的制式必然要用尖头弹。7.92mm圆头弹和7.92mm尖头弹直径不一样 根本无法通用 其实和增加一种口径没有什么区别。7.92mm圆头弹的枪口动能在3000J左右 后坐力的问题并不突出 所以民国初年采用7.92mm圆头弹是符合中国国情的。但如果换成7.92mm尖头弹 枪口动能达3800J 后坐力过大的问题就显现出来了。7.92mm尖头弹既不能简化后勤 又不适于中国士兵的体质 显然不是一种好的选择。反正也是要增加一种口径 为何不干脆采用更适合中国战场的枪弹呢？（4）备选方案如果不追求步枪和机枪弹药统一 则步枪弹用6.5×50mm有坂弹 机枪弹用7.92×57mm毛瑟弹（尖头） 完全能发挥各自的长处。况且这两种子弹国内的生产经验都比较丰富 生产线是现成的 投入资源较少 大批量生产很容易。（二）步枪抗战前 各路军阀从各种渠道进口了大量步枪 种类五花八门 国内各个兵工厂也仿制了多种步枪。归结起来看 进口步枪中 以德国毛瑟98系列和日本三八式数量较多。其次是奥匈曼利夏M1895、意大利卡尔卡诺M1891和苏俄莫辛-纳甘 前两者都是一战后的作为剩余武器出口到中国；后者一部分是苏俄内战后流入中国 另一部分则是苏俄在国共合作北伐时期的军援。其他种类的步枪比如英国李恩菲尔德、法国勒贝尔1886等进口数量都较少。而美国斯普林菲尔德M1903和M1917是在抗战后期才作为军援进入中国的 早期国内并没有装备美制步枪。国内自行制造的仿制品中 主要是汉阳造、毛瑟98系列和三八式。（1）30年代各种步枪的优缺点分析上述众多列举的步枪中 按技术和性能来讲 有的已经过时 不太适合二战的环境。法国勒贝尔1886是世界上第一种使用无烟火药的枪械 年代最老 性能最差。汉阳造源自德国1888式委员会步枪（注意不是毛瑟） 经过了中国人的改进 国内制造和使用的经验都比较丰富 有利于扩大产量 简化后勤；然而其性能已经落后于时代 大规模装备只能是浪费资源。奥匈曼利夏M1895和意大利卡尔卡诺M1891性能相对好一些 但也比较过时。而几大军事大国的制式步枪 苏俄莫辛-纳甘、英国李恩菲尔德、德国毛瑟98、美国斯普林菲尔德M1903和日本三八式步枪各有特色 性能差别不是很大 作为手动步枪都能满足二战的环境。当然 和半自动步枪、冲锋枪没有可比性 战术要求不一样。莫辛-纳甘易于制造 维护简单 但枪机设计较为复杂 操作感觉有些笨拙 人机功效较差。日本三八式射击稳定 后坐力小 但杀伤力的确弱一些。李恩菲尔德在手动步枪中弹容量最大 射速最快。总体而言 德国毛瑟98和美国斯普林菲尔德M1903的精度、杀伤力、工艺性、可靠性等指标比较平衡 综合性能在上述所有步枪中最好。其实美国斯普林菲尔德M1903本来就是德国毛瑟98的美国版仿制品 只不过改了口径而已 两者性能类似。 抗战前制式步枪的选择 一是要考虑步枪的性能 不一定最好 但也不能过时；二则要考虑本国的兵工现状 最好是选择有仿制经验的 有利于扩大产量。当然 仅限于手动步枪 半自动步枪根本还没有成熟 也不是中国能玩得起的。三八式步枪以阎锡山的太原兵工厂仿造较多 其他兵工厂如广东兵工厂、巩县兵工厂等主要仿造的都是毛瑟98系列。其他诸多步枪几乎都没有仿制经验 如果另起炉灶需要时间 不能满足国军急切的装备需求。在保证性能不落后的前提下 自然要选择对兵工设备工艺调整量最小 对后勤供应体系变化最小的步枪 所以制式步枪选择毛瑟98系列中的一种是最佳方案。国民政府的大方向是正确的 但在具体选型上却出了偏差。（2）长枪管和短枪管的差异毛瑟98系列在欧洲有G98（最初型号）、98a、98b、1924标准型、FN 1930和98K等 国内仿制品有元年式、四年式、辽十三式、巩造98式和中正式等。按枪管的长短又可分为长枪管和短枪管两大类 G98、98b、元年式、四年式、辽十三式、巩造98式均为长枪管；98a、1924标准型、FN 1930、98K、中正式则为短枪管。三八式步枪则是典型的长枪管。相对而言 长管步枪的年代早一些 枪管长度在750mm左右；短管步枪的年代晚一些；枪管长度在600mm左右的步枪。短管步枪是进入二十世纪后的战争形式变化和技术发展的产物。在第一次世界大战之前 陆战的主要形式是野战环境之下的大规模运动战。比较长的步枪有利于士兵在开阔地上击中距离更远的敌人 在白刃拼刺时也具有显而易见的优势 因此各国步兵装备的步枪普遍比较长。到了一战时期 阵地战取代野战成为主流的陆战形式。长管步枪拥有750mm的枪管和最大射程远至2km之外的表尺 虽然在理论上可以击中极远距离的目标 但是在这个距离上击中在战壕中只露出头和手臂的敌人的概率极小。同时较长的枪身也造成了在战壕里活动不太方便。同时 进入二十世纪二三十年代后 随着技术的发展 发达国家军队机械化程度日益提升。重武器和装甲车辆的装备数量的增加强化了远距离火力打击能力 步兵交战的距离则缩短到不超过400m 不再需要靠长枪管来保证远距离的精确射击。同时乘车作战的模式也开始普遍 较长的枪身不便于随车携带。基于上述的两个原因 较长的枪身变得弊大于利。因此各国纷纷将原来的长管步枪换成了短管步枪。抗战前 国民政府最终选择了短管步枪 即基于1924标准型的中正式步枪作为国军的制式步枪。从表面看 似乎是跟上了发达国家步枪更新的潮流 但仔细研究之下 事实却并非如此。问题的根源还是在当时中国的工业水平 无法提供足够的重武器以保证远距离火力打击 弹药补给能力也非常薄弱 无法保证火力的持续性 机械化更是空谈。所以中国战场的陆战形式事实上还停留在一战之前的水平上 总体上双方决定胜负的仍然是步兵集群在野战战场上的对决。这种客观环境决定了长管步枪才更符合中国战场的需求：一是瞄准基线长 射击精确度高；二是枪管长使火药燃烧充分 降低了枪口焰 提高了士兵隐蔽和生存能力；三是有利于白刃战。国民政府和国军的相关负责人没有仔细考量当时中国的工业水平 高估了国军炮兵和装甲兵发展速度 高估了国军的弹药补给能力 对于白刃战在迫在眉睫的中日战争的作用认识不足 因此超前地采用了中正式步枪作为制式步枪。中正式步枪由于枪身短 拼刺能力较弱 于是不得不配备了很长的刺刀。即便如此 中正式安上刺刀后仍然比安了刺刀的三八式短一截；而刺刀太长外加制造工艺不过关 又极易变形和损坏。结果是既在火力上处于劣势 又在白刃战也处于劣势。（3）长枪管毛瑟步枪适合中国战场的需要通过上述的分析可以看到 抗战时期中国军队采用长管步枪才是符合国情的选择。在当时国内已经有的长枪管毛瑟98系列仿制品中 有元年式、四年式、辽十三式、巩造98式。元年式和四年式同出一脉 是民国初年的仿制品 元年式最初采用6.8mm口径 后来改为7.92mm口径就变成了四年式 两者都使用圆头弹 规格较老。辽十三式量产于1924年 为奉天兵工厂所造 和国内其他毛瑟步枪仿制品有所不同 可以说是毛瑟和三八式的混合体。巩造98式量产于1933年 为巩县兵工厂所造 是在G98的基础上参照辽十三式的图纸改进而来 采用尖头弹 规格相对较新。综合比较下来 以巩造98式为基础 并且在口径上做改进 使用7×57mm毛瑟步枪弹 成为一支全新的制式步枪（姑且称之为巩造新98式）。这样 从子弹杀伤力看 新枪要超过三八式；从使用角度来看 新枪的后坐力较小 便于精确射击和士兵训练；从白刃拼刺能力看 新枪不次于三八式。在中国军队应该以巩造98式为基础 缺乏重武器的情况下 该新枪作为中国士兵手中最基本的轻武器 性能超过了日军 将成为抗战的有利保障。（4）备选方案对应步枪弹的备选方案 如果步枪弹用的6.5×50mm有坂弹 则制式步枪干脆就用三八式。实际上 三八式是一支不错的步枪 绝不是某些无脑写手笔下的废物。该枪除了枪身长 后坐力小带来的好处 还有一些独创之处。比如它的防尘盖 不仅是该枪的标志性符号 也是该枪最大的亮点。安装防尘盖 能够有效地阻止泥沙、灰尘进入枪机 减少了在尘土飞扬的战场上发生故障的概率 很有实战价值 也使全枪的外观显得干净利落。安装这么一个盖子 工艺要求并不复杂 生产成本也并不昂贵 可谓是以小的代价完成了大的贡献。其它比如它的枪机、保险机、瞄准装置、枪托 都有其特点。所以除了杀伤力稍弱一些 三八式其实还是很适合在中国战场使用的 国内也有丰富的仿造经验 可以作为备选制式步枪。（三）机枪机枪是步兵最基本的火力支援武器。最初的机枪都是重机枪 轻机枪出现于第一次世界大战前后 通用机枪则要到在20世纪30年代才被德国首先装备。民国时期各路军阀最初装备的机枪都是重机枪；轻机枪起初数量很少 直到20世纪20年代后期才开始大量装备；通用机枪更是在1949年前都不曾出现在中国。网上的军事玄幻小说中 动不动拿MG34、MG42装备国军 根本不考虑当时的中国是否造得出、玩得起这种武器。MG34的确先进 但工艺复杂 以中国当时的工业水平 制造难度极大 比如为保障高射速所需的金属弹链就造不出来。所以在机枪的选择上 不能好高骛远 还是老老实实按照重机枪和轻机枪分别装备。1. 重机枪重机枪最初由英籍美国人马克沁发明。重机枪可分为两类 水冷式和气冷式 在30年代之前 世界上的重机枪主要分为三大体系。德国马克沁MG08 苏俄马克西姆M1910 英国维克斯都是从马克沁机枪发展而来 为水冷式。法国哈奇开斯重机枪开了气冷式重机枪的先河 日本的明治三十八年式 大正三年式都仿自哈奇开斯。美国则采用勃朗宁式重机枪 M1917为水冷式 M1919为气冷式。历史上的中国主要仿制了其中两种 仿德国马克沁MG08的民二四式和仿美国勃朗宁M1917的三十节 其他类型都比较少。到了30年代中后期及二战期间 新出现的捷克ZB-53 意大利布雷达M37 日本九二式 苏俄郭留诺夫SG-43等重机枪 都是气冷式 反映了气冷式取代水冷式的趋势。水冷式重机枪只要水没有蒸发完 就能维持枪管的温度不超过100度 所以持续射击能力强 对枪管钢材和加工的要求较低。缺点是重量较大 移动不方便；射击过程中会蒸发水汽 容易暴露位置；一旦缺水或水筒被打坏 就无法使用。气冷式在射击过程中会没有水汽产生 不容易暴露位置；使用不受水的限制。缺点是枪管升温快 需要经常停顿冷却或更换枪管 持续射击能力差 对枪管钢材和加工的要求较高。最初的气冷式重机枪如法国哈奇开斯 日本明治三十八年式的重量和水冷式差不多 因此优势不明显。但后来出现的美国勃朗宁M1919A4 捷克ZB-53 意大利布雷达M37 苏俄郭留诺夫SG-43的重量都大为减轻 逐步取代了本国的水冷式重机枪。原因在于现代战争的火力打击能力增强 重机枪长时间保持在一个阵地容易被迫击炮、无后坐力炮等火力消灭；重型武器的增加降低了部队对重机枪的依赖；战术的进步也要求机枪火力能伴随步兵行进。其持续射击能力强的优点变得多余 而其重量较大 移动不方便 受水限制的缺点凸显出来。所以气冷式取代水冷式是大势所趋 后来的通用机枪则完全是气冷式的天下了。虽然世界趋势如此 但中国的情况却有其特殊性。第一 30年代之前 中国的冶金工业极为薄弱 难以保证气冷式重机枪对钢材和工艺的要求；第二 由于缺乏重型武器和机枪数量不足 战斗中非常需要重机枪能持续射击提供火力支援。所以在中国战场 至少是抗战前期 水冷式更符合兵工生产和实战的需要。因此在30年代 仿制德国马克沁MG08的确是重机枪的最优选择。当然 最好是把口径改成7mm 使用前面说的7×57mm毛瑟步枪弹 做到步机枪弹药统一。当然 到了抗战后期 可以考虑仿制气冷式重机枪 比如美国勃朗宁M1919A4或苏俄郭留诺夫SG-43 也可以研究把马克沁改成气冷式。（这是可行的 历史上联勤部二十一兵工厂1945年开始研究将水冷式马克沁改成气冷式 于1947年成功造出样枪）。2. 轻机枪世界上最早的轻机枪是1905年问世的丹麦麦德森轻机枪。由于轻机枪重量轻 能伴随步兵快速机动 因此第一次世界大战开始大量装备各国军队。中国很早就进口并仿制过轻机枪 如丹麦麦德森、法国哈奇开斯M1909、法国绍沙M1915、日本大正十一年式（就是歪把子） 但这些轻机枪年代较早 性能不佳 因此装备和仿制数量都很少 不成规模。直到20世纪20年代后期 中国才开始大量装备并仿制轻机枪。仿制品最多的是捷克ZB26（著名的捷克式） 其次为瑞士启拉利。抗战前进口但没有仿制过的有法国哈奇开斯M1922、比利时勃朗宁FN1930、芬兰拉提M26和德国MG13。抗战中进口或援助的有苏俄捷格加廖夫DP、美国勃朗宁M1918和加拿大勃然式。除去早期的轻机枪 上面列举的轻机枪中 除了加拿大勃然式 在30年代前期都已经面世。大部分轻机枪有其优点 但缺点也比较明显 比如 瑞士启拉利结构最简单 制造最容易 但精度较差；芬兰拉提M26精度很好 但零件太精密 加工难度较大；捷格加廖夫DP弹容量较多 但弹盘的故障率较高 全枪重量和尺寸都偏大 携带不变 等等。而捷克ZB26和比利时勃朗宁FN1930的精度、杀伤力、工艺性、可靠性等指标比较平衡 综合性能更好。捷克ZB26和比利时勃朗宁FN1930相比有个优势 就是能够快速更换枪管 这是一个里程碑式的创造。气冷式重机枪可以通过采用重枪管加大热容量 开散热孔的方式来延缓升温 而轻机枪为了控制重量很难采用重枪管。射击一段时间后枪管发烫 就必须停下来等待冷却 否则不但子弹失去准确性 还会影响枪管寿命。能够快速更换枪管 就可以保持火力的连续性 在战场上好处是巨大的。捷克ZB26开创了先河 在其之后的轻机枪纷纷添加了该项功能。再加上捷克式结构简单 容易操作 历史上中国军队选择捷克式作为制式轻机枪应该说是个明智的选择。然而捷克式也有一个不足之处 就是弹匣置于枪身上方。这带来两个问题 一是其瞄准装置只能采用偏出枪体的瞄准方式 虽然并不影响射击的精确性 但是影响了射手的视线；二是整支枪的重心相对偏高 造成枪容易倾斜 转动射击左右方向时也不好控制枪身。而比利时勃朗宁FN1930的弹匣在枪身下方 就没有这两个问题。那么 有没有一种轻机枪 结合了捷克ZB26和比利时勃朗宁FN1930两者的优点呢？有的 那就是比利时勃朗宁FN D型 它是勃朗宁系列中的最新、最先进的改进型 定型于1932年 具备快速更换枪管的能力。（“D”这个字母来自法语“Demontable”——意思是“可拆卸”。）它的基本弹匣容量和ZB26一样为20发 有些偏少 但是弹匣在枪身下方 所以还有改用大容量弹匣或者弹鼓的潜力。比利时勃朗宁FN D型的各项指标都很出色 综合性能一流 制造也不比捷克式复杂 非常适合当时的中国。而且中国是在20世纪20年代后期才仿制捷克式 还没有形成大规模 选择一种新型号并不会影响原有的兵工生产和后勤保障体系。中国军队应该选择比利时勃朗宁FN D型作为制式轻机枪 并和重机枪一样 把口径改成7mm 使用7×57mm毛瑟步枪弹 做到步机枪弹药统一。3. 备选方案备选方案就很简单 和历史上的做法一样 直接使用马克沁水冷式重机枪和捷克ZB26式轻机枪 它们的优缺点在前面已经叙述过 不再重复。轻重机枪的口径都不需要更改 直接用7.92×57mm毛瑟弹。虽然捷克式轻机枪不如比利时勃朗宁FN D型 但胜在仿制经验丰富一些 对工业生产能力的要求低。（四）手枪和冲锋枪1. 手枪民国前期中国进口的手枪五花八门 品种繁多 仿制也不少。总体来说分为三大类 一类是左轮枪；一类是大名鼎鼎的毛瑟军用手枪 俗称盒子炮；剩下的就是各种半自动手枪 俗称“撸子”。其中左轮枪问世年代最早 明显已经不适合现代战争 不用考虑。中国在20世纪前半期最流行的手枪莫过于盒子炮 诞生于1896年的德国毛瑟兵工厂 历史上中国曾大量进口并仿制。盒子炮在出生地欧洲并不受重视 没有一个国家把它列为制式武器。因为它结构复杂 价格比一般的手枪高几倍 重量和尺寸也大；和步枪冲锋枪相比威力又过小；显得高不成低不就。它在中国的流行其实是因为民国初年连年内战 国际联盟对中国实行了长达十年的“武器禁运” 步枪和冲锋枪都不能合法地进口 而各类手枪却不在受禁之列 可以堂而皇之地大量进口。盒子炮的枪管长 弹容量大 因此射程、精度和火力持续性都超过了普通手枪 能适应多种场合。它在中国其实是作为冲锋枪的简化版替代品来使用 以补充中国各路军阀步枪冲锋枪数量的不足。民国初年的军阀战争烈度都不大 盒子炮恰好能发挥其长处 风骚一时。但替代品就是替代品 各方面的性能毕竟不能和正规的冲锋枪相提并论。到了抗日战场 正面战场的战争烈度大大增强 盒子炮这种替代品是不能满足战术需要的 近战火力还是应该以正规的冲锋枪为主。历史上 无论是国共双方的军队 随着冲锋枪数量的增加 盒子炮逐渐被淘汰就是无可争议的事实。与其生产盒子炮 还不如把有限的资源用于多生产一些冲锋枪。当然 在敌后的游击战中 盒子炮还是能发挥很大作用的。手枪的选择 则应真正回到其自卫武器的定位。在民国早年的各种半自动手枪中 以勃朗宁系列手枪最受青睐 有“一枪二马三花口”的说法 指的是M1900（枪牌撸子）、M1903（马牌撸子）、M1910（花口撸子）。不过这是指它们问世的时间顺序 而不是性能排列。从性能看 以M1903最佳 M1910次之 M1900最差。这些早期的勃朗宁手枪发射的子弹威力不足 弹容量也小 只能用于自卫 在其它战术领域如侦察 渗透等方面的使用则有缺陷 多用性差一些。后来的勃朗宁M1911采用0.45英寸（11.43mm）柯尔特手枪弹 威力强大 停止作用好 美军特种部队至今仍在使用 但它的后坐力较大 不适合中国人的体格。最后出现的勃朗宁M1935式手枪 采用9mm帕拉贝鲁姆手枪弹 弹容量大 达到13发 性能也极为出色 后坐力适中。总体来看 勃朗宁M1935式手枪是制式手枪的最佳选择。2. 冲锋枪冲锋枪诞生于一战 但在一战到二战之间的这个时期发展缓慢。大量优秀的冲锋枪是在30年代末和二战期间诞生的 比如德国MP 38/40、意大利伯莱塔M38、英国斯登、苏俄波波沙、美国M3等。在30年代前期 可选择仿制的冲锋种类不多 无非是德国MP18、美国汤姆森和芬兰索米。其中性能以芬兰索米最佳 但其加工过于精密 仿制难度和成本较高；美国汤姆森重量偏大 结构复杂 同样不利于大量生产；只有德国MP18 结构简单 操作方便 适合中国这样工业基础薄弱的国家。MP18伯格曼冲锋枪 由于枪管上有多空散热套 在中国被形象地称为“花机关”。它只有30几个零件 零件也并不精密 不需要高精度的加工工具 即使零件出现少许误差 也不会影响射击的精度和稳定性。历史上 中国不少兵工厂如上海、金陵、广东、巩县等都曾经仿制过 可见其结构之简单 工艺之普通。MP18的性能相当不错 坚固耐用 射击精度较好 易于操作和维护。在一战中 MP18参战不过几个月 就取得了很好的战果。在德军投降以后 英法立即下令 德军未来都不得继续研究和装备MP18冲锋枪 可见其对英法军队打击之大。因此中国应采用MP18冲锋枪作为制式冲锋枪 加强近战火力和战术灵活性。3. 手枪弹大多数国家的手枪和冲锋枪用同一种子弹。20世纪30年代世界上比较流行的手枪弹主要有：9mm帕拉贝鲁姆手枪弹 7.65/9mm勃朗宁手枪弹 0.45英寸（11.43mm）柯尔特手枪弹 7.63mm毛瑟手枪弹。9mm帕拉贝鲁姆手枪弹尺寸适中 威力大 精度佳 停止作用好。勃朗宁手枪弹的优点是精度好 后坐力小 容易控制 缺点是军用威力不足。0.45英寸柯尔特手枪弹的优点是威力最大 停止作用最好 缺点是后坐力大 不容易控制 子弹体积也大 携弹量少。7.63mm毛瑟手枪弹的优点是初速高 射程远 侵彻力强 精度良好 缺点是弹头口径小 质量小 近距离容易穿透 停止作用差。从现代的眼光看 0.45英寸柯尔特手枪弹威力最大 停止作用最好 9mm帕拉贝鲁姆手枪弹性能最平衡。所以帕拉贝鲁姆弹和柯尔特弹在21世纪继续流行 尤其是帕拉贝鲁姆弹已成为世界通用标准弹 使用最广泛 装备数量最多。而另外两种手枪弹则已经逐渐消失 是有道理的。在中国 大部分盒子炮和部分的MP18伯格曼冲锋枪都使用7.63mm毛瑟手枪弹 这是中国使用量最多的手枪弹。勃朗宁M1935手枪 小部分盒子炮和部分MP18伯格曼冲锋枪使用9mm帕拉贝鲁姆手枪弹。勃朗宁M1903和M1910使用的是7.65mm或9mm勃朗宁手枪弹。勃朗宁M1911手枪和汤姆森冲锋枪使用0.45英寸（11.43mm）柯尔特手枪弹。根据上面对各种手枪弹的性能分析 再考虑到已经选定勃朗宁M1935手枪和MP18伯格曼冲锋枪作为制式手枪和冲锋枪 那么抗战前的中国以选择9mm帕拉贝鲁姆手枪弹作为制式手枪弹就顺理成章了。4. 备选方案手枪方面 分为战斗手枪和自卫手枪两种制式。考虑到毛瑟军用手枪在中国的使用和仿制经验都比较丰富 直接作为战斗手枪 配备基层军官、警卫人员、侦察分队和二线战斗人员等。中高级军官则另外配备合适的自卫手枪 在民国前期的自卫手枪中 以发射9mm勃朗宁手枪弹的M1903（马牌撸子）性能最佳。好在中高级军官配枪数量很少 增加一种制式对后勤的影响可以忽略。备选方案的冲锋枪制式不变 仍是MP18伯格曼。但是枪弹使用7.63mm毛瑟手枪弹 和盒子炮保持一致。（五）轻型火炮（迫击炮和山炮）1. 迫击炮迫击炮自问世以来 一直是支援和伴随步兵作战的一种有效的压制兵器。它的射角大 弹道弯曲 特别适合于用来对付遮蔽物后方的目标；操作简单 装弹容易 射速很高（20～30发/分） 火力猛；质量轻 体积小 中小口径迫击炮可以人背马驮 打了就跑 能快速转移阵地 机动性强。 对于当时缺乏重武器的中国军队来说 迫击炮是一种非常实用的武器。最为关键的是 迫击炮的技术难度和成本都比其他火炮低得多 易于大规模生产。一般火炮身管要承受很大的膛压 需要高品质的钢材 加工要求也很高 这对30年代的中国工业水平是个很大的障碍 难以大规模制造。迫击炮则不同 由于膛压低 只需要普通的无缝钢管就可以制造 非常适合中国国情 可以迅速扩大产量。历史上 中国早在20年代就有仿制迫击炮的经验 但在抗战前对迫击炮的战术作用认识不足 制造和装备数量并不多。开战后吃了日军掷弹筒不少亏后 才加大了迫击炮的产量。如果能够早日仿制比较先进的迫击炮 并大量装备 必将取得良好的效果。30年代最为出色的迫击炮莫过于法国布兰德60mm和81mm迫击炮 中国应当以此为基础 发展60mm、82mm、120mm三个级别的口径。在抗战之初 60mm小口径装备到营 82mm中口径装备装备到团 120mm大口径装备到师 形成梯次火力。随着产量的扩大 可以考虑把60mm口径装备到连 82mm装备到营 120mm装备到团 逐级下放 进一步增强步兵伴随火力。2. 山炮山炮其实是轻型榴弹炮 它通常可以分解后由马驮载 或者直接由马拖拽 特别适合山地作战 因此才冠名为山炮。20世纪30年代 世界主流山炮一般都为75mm口径 重量都在1000kg之内。山炮的技术难度不算高 中国从清末开始就有山炮的仿制经验。清末江南制造局于1905年仿制德国克虏伯14倍径75mm山炮 称沪造克式75mm山炮。汉阳兵工厂于1921年 太原兵工厂于1924年 奉天兵工厂于1925年 分别仿制日本四一式75mm山炮成功 称汉10年式、晋13年式、辽14年式75mm山炮 其中以太原兵工厂产量最大。可见 国内的兵工企业有制造山炮的能力。因此在进口先进山炮的同时 也要积极加以仿制 争取早日实现国产化。历史上 中国进口了一批瑞典博福斯M1930式75mm山炮 属于当时世界上最先进的山炮之列 重量约700多kg 射程超过9km 精度极佳。相比之下 国内仿制量最大的日本四一式山炮设计年代较早 虽然重量较轻 不到600kg 但射程也较短 约6km多 总体性能不如博福斯山炮。和博福斯山炮性能相近的其他75mm山炮有法国施耐德M1923式、捷克斯柯达M1928式和美国M1A1（又称M116）。一战之后 为了规避《凡尔赛条约》的限制 德国把一些军事工业转移到邻国去发展 德国克虏伯军火工业就收购了瑞典博福斯兵工厂部分股权 并开展合作研究。在中德军事合作的前提下 取得博福斯山炮的技术相对于其他国家可能性大一些。因此采用博福斯M1930式75mm山炮作为制式山炮是最佳选择。3. 其它支援火力掷弹筒和九二式步兵炮是日军特有的武器 曾经在中国战场发挥了很大的作用。但是它们退出历史舞台的速度又很快 二战后就再也没有其它国家使用过类似武器。从性能上说 它们都不如迫击炮 它们的作用只限于特定的历史条件和特定的战场 也和日军最初对迫击炮不重视有关。从原理上来说 掷弹筒就是一门超轻型的迫击炮。它的优点是重量很轻 可以单兵携带 隐蔽性很。它的缺点一是没有迫击炮的瞄准具 精度不足 所以必须经过长时间训练才能掌握好使用技能；二是杀伤力和射程也远不如60mm口径的迫击炮。日军可以提供足够的时间和资源给士兵来训练使用这种单兵武器 中国却没有这个条件。有限的兵工资源只能优先满足更有效的武器 除了小口径迫击炮 还应该生产枪榴弹筒来加强一线步兵的支援火力。枪榴弹筒杀伤力和掷弹筒相似 但可以依托步枪来瞄准和发射 精度相对较高 训练也更简单。二战后 掷弹筒迅速淘汰 枪榴弹筒却逐渐演化为枪榴弹发射器 继续装备一线步兵 就很能说明两者谁更有生命力。步兵炮诞生于一战 二战后就趋于消亡 生命周期十分短暂。这种武器的最大特点在于能同时曲射和直射 但两方面的性能都比较平庸。以日军九二式步兵炮为例 口径为70mm 重量却达200kg；80mm级别的迫击炮威力射程和它差不多 射速更快 重量却只有60kg左右 而结构更是简单多了。造一门九二步兵炮的资源投入完全能够造好几门82mm迫击炮 所以用于曲射武器 中口径迫击炮远胜过步兵炮。步兵炮超过迫击炮的地方在于它的直瞄射击能力。但由于炮弹初速太低 才200m/s 进攻作战中只能对付轻型野战工事 也就是木土工事和较薄弱的砖石工事 真正的钢筋混凝土工事 它是打不掉的；防御战中 反装甲能力则更弱。直射武器 与其使用步兵炮 不如多装备一些反坦克炮 无论在进攻还是防御战中 能起的作用更大。总体看来 步兵炮的曲射费效比不如迫击炮 直射费效比不如反坦克炮。九二步兵炮在中国战场大放异彩大紫 只因为中国军队的迫击炮和反坦克炮数量实在太少 没有办法压制它；而到了太平洋战场 在美军的迫击炮和反坦克炮群面前 根本没有用武之地。反过来对于国军来说 在资源有限的情况下 更应该优先装备迫击炮和反坦克炮。综上所述 掷弹筒和步兵炮都不适合作为国军的制式武器 枪榴弹筒则应该作为一种制式武器装备一线步兵。（六）重型火炮（野炮和榴弹炮）重型火炮的远程火力打击对现代战争的重要性是毋庸置疑的。不过在20世纪30年代 中国的“重炮”和欧洲战场的“重炮”概念完全不同。欧洲师一级的标准支援火炮大多是75mm野炮和105mm（或100mm）榴弹炮 比如比利时、罗马尼亚军队；德国、法国等军事强国的精锐部队则是105mm榴弹炮和150mm（或155mm）榴弹炮。日本陆军在抗战初期 一个师团的炮兵联队或是装备36门75mm山炮和75mm野炮（驮马制） 或是装备36门75mm野炮和120mm榴弹炮野炮（挽马制） 火力比欧洲陆军要差一些。无论是欧洲还是日本 105mm及以上级别的加农炮、150mm及以上级别的榴弹炮才算是重炮 一般都编组成独立的重炮部队。而对重武器缺乏的中国军队来说 75mm以上口径的野炮、榴弹炮就已经算是“重炮”了。抗日战争的烈度虽然和欧洲战场相比远远不如 但一定程度的重炮支援还是很有必要的。博福斯75mm山炮的性能虽然优秀 但9km的射程毕竟有限 是无法承担远距离火力支援任务的 中国战场的重炮至少也要保证10km以上的射程。20世纪30年代有好几种比较优秀的150~155mm口径的榴弹炮问世 包括德国莱茵金属s. FH 18式 捷克斯柯达M1934式 瑞典博福斯M31式 日本九六式等。前三者性能类似 重量都达到5吨以上；日本九六式的重量稍轻 为4吨多 但射程也近一些。历史上国民政府在德国顾问的建议下 采购了48门s. FH 18式150mm榴弹炮 编成两个炮兵团。它们的威力大、精度好 在抗战中发挥了一定的作用。但是客观地说 150mm口径的重炮并不适合当时的中国战场环境。这个重量级别的火炮通常需要用汽车拖拽 用马拉的效率很低。在欧洲 依托发达的公路网 可以方便地实现机动。但20世纪30年代的中国 道路状况非常差 特别是山区和水网地带 可供汽车行驶的道路极少 重炮机动受到极大的限制。同时 中国空军的实力处于绝对弱势 战场的制空权将迅速丧失 炮兵一旦开火 就会处于日军航空兵打击的威胁之下 转移阵地不便大大降低了重炮的生存性。因此 s. FH 18式150mm榴弹炮在中国实际发挥的作用远没有预想的大 很多情况是需要火力支援的地方去不了 到了地方也不敢随时开炮。更何况150mm榴弹炮的价格极为昂贵 性价比并不高。所以 中国的“重炮”首先要考虑的就是便于机动 重量不宜超过2吨。这样在路况较好时就用汽车拖拽 路况不佳时用马拉也很方便 机动性大大提高 既能扩大火炮的使用地域 也增强了火炮的生存能力。历史上淞沪会战后期国军撤退时 由于一座公路桥被工兵布雷 炮10团的汽车无法通过 不得已只能把部分150mm榴弹炮推入河中抛弃。如果是2吨以内的火炮 也许就能选择小路用马拉过河 或者用船运过河 避免装备损失。考察当时先进火炮的技术指标 抗战前的中国应选择75mm口径（或接近）的野炮和105mm口径（或接近）的榴弹炮 才能同时满足重量2吨内和射程10km以上的要求。而且价格肯定比150mm榴弹炮便宜 同样的预算可以多买一些。这些重炮应以团为单位 编组成独立的预备炮兵部队 由战区一级的指挥部掌握 根据需要加强到重点战场提供火力支援。75mm野炮射速较高 105mm榴弹炮炮弹威力较大 两者配合使用相得益彰。在具体型号方面 应选择德国le. FK 16式75mm野炮和le. FH 18式105mm榴弹炮 前者重量约1.5吨 后者重量约1.9吨 两者射程都超过10km 达到了12km左右。优先选择德国的火炮是考虑了30年代中德军事合作的背景 可以取得贷款并以矿产还贷 比较优惠。其他国家也有性能类似的火炮 比如法国施耐德M1927式85mm野炮和M1934式105mm榴弹炮 捷克斯柯达vz30系列的76.5mm野炮和100mm榴弹炮等。但这些火炮都需要现款支付 财政负担较大 不如德国炮经济。进口75mm野炮和105mm榴弹炮对中国的兵工生产也有积极的作用。因为它们的仿制难度比150mm榴弹炮小得多 炮弹制造难度也比150mm炮弹容易 能够从一个较低的起点出发 逐步提升 以减少对进口的依赖程度。le. FK 16式75mm野炮和le. FH 18式105mm榴弹炮对抗日军各师团的队属炮兵绰绰有余 但比日军的独立重炮部队装备的新式大口径榴弹炮和加农炮还有不小的差距。尤其是日军的加农炮 如92式105mm加农炮和89式150mm加农炮 96式150mm重加农炮等 性能都很优秀 射程远远超过s. FH 18式150mm榴弹炮。这是当年的中国军队怎么也无法抗衡的先进武器。所以中国军队必须放弃和日军新式火炮的正面对抗 把预备炮兵的作用定位在能够压制日军师团队属炮兵就行了。好在日军新式火炮数量并不多 而且重量都比较大 受道路条件限制 转移阵地比较费时。完全可以利用le. FK 16式和le. FH 18式实施打了就跑的机动战术 制造重点战场的局部优势 取得良好的战果。（七）反坦克和防空武器在抗战中 日军的飞机和坦克对于中国军队的威胁非常之大。尤其是在战争初期 作战地域处于中国东部平原地带 对日军的飞机和坦克发挥作用有利。建设一支强有力的空军和装甲部队需要长期而且巨大的投入 包括装备采购 人员培训 机场建设 后勤保障等等。以当时中国的国力而言 想在短期内建立全面超过日本的空军和装甲部队是力不从心的 只能维持少数精干的空军和装甲部队 用于一些重点战场。形势决定了中国军队对日军的飞机和坦克将长期处于防御状态。因此 引进一批有效的防空和反坦克武器 不失为成本比较低廉 见效比较快的对抗手段。1. 反坦克炮日军的坦克都不重 普遍装甲薄弱 所以一般37mm以上的反坦克炮都能对付。考察30年代前期的反坦克炮 可选择的反坦克炮有德国Pak36式37mm反坦克炮 瑞典博福斯37mm反坦克炮 捷克斯柯达vz34式37mm反坦克炮 比利时M1931式47mm反坦克炮 奥地利百禄B?hler 式47mm反坦克炮。这些炮的性能相差不是很大。威力以比利时的47mm反坦克炮最大 但重量也最重 超过500kg。其它炮都在450kg以下。 奥地利百禄B?hler式47mm反坦克炮的重量很轻 不超过350kg左右 机动性极好。它最大的特点是射角很高 其它反坦克炮的仰角只有约20度 它的仰角则达到近60度。这样高的仰角使得百禄式反坦克炮可以作为轻型山炮提供火力支援 比一般的反坦克炮用途更广。而且47mm的口径可以发射比37mm口径重一倍的炮弹 杀伤力更有保证。意大利的布雷达M1935式47mm反坦克炮其实就是百禄式 是从奥地利取得了许可证后生产的。意大利军队就把它同时用作反坦克炮和轻型山炮。对于缺乏武器的中国军队来说 有这样一种轻便而多用途的火炮实在是很经济的选择。2. 反坦克枪受限于财政状况 国军不可能采购大量的反坦克炮 所以需要更廉价的反坦克枪作为补充 装备一线步兵。30年代前期世界上的反坦克枪种类不多 只有德国毛瑟M1918式13.2mm反坦克枪和索罗通S18-100式20mm反坦克枪可以选择。其它在二战中有名的德国Pzb38反坦克枪 英国博伊斯反坦克枪 苏联PTRD 1941反坦克枪等都要在30年代末才出现。从威力看 自然是索罗通S18-100式20mm反坦克枪更强 但是它的重量达到40多千克 不太适合中国士兵。德国毛瑟M1918式13.2mm反坦克枪不到20千克 价格更便宜 虽然穿甲能力差一些 但对日军的薄皮坦克还是很有效果的。反坦克枪的威力远胜一般步枪 除了装甲目标外 也可以用来对付工事 车辆 火力点等目标。现代的反器材步枪就是从反坦克枪发展而来。3. 高射炮应该说 国民政府对防空作战是有一定的认识和准备的 也进口了一批高射炮 包括20mm小口径机关炮 和瑞典75mm、德国88mm的大口径高射炮。这种组合缺乏针对性 费效比不太高。防空作战分为要地防空和野战防空。一般而言 大口径的高射炮重量大 射速慢 多为手动装填 射程远 针对高空目标 执行要地防空任务；中小口径的高射炮重量轻 射速快 多为自动装填 射程近 针对中低空目标 执行野战防空任务。在欧洲战场 飞机种类齐全 尤其是英美装备了大量战略轰炸机 因此大中小口径的高射炮都有必要装备 形成覆盖整个空域的火网。而对国军来说 则不宜装备大口径高射炮。第一 在中国战场 日本陆海军航空兵的飞机虽然比中国先进 却比欧美强国落后许多 大型轰炸机很少 只有部分中型轰炸机 大部分是轻型的战斗机和攻击机。针对日军航空兵 大口径高射炮从技术角度来说性能显得浪费。第二 大口径高射炮价格昂贵 采购数量过少又不足以形成火网 战术效果打了折扣。第三 大口径高射炮重量比较大 移动不便 比如德国88mm高炮重达5吨 只能固定阵地 武器的利用率不高。因此国军应该以中口径的高射炮为主 辅以小口径的高射炮。在二战中 性能最好的中口径高射炮无疑是瑞典博福斯40mm高射炮。无论是同盟国还是轴心国 都大量制造 广泛使用 将其视为标准防空武器。它的精度好 可靠性高；威力和射高均优于20mm轻型高炮 射速又高于75mm以上的重型高炮 能够有效对付中低空的目标；同时重量不超过2吨 具有较强的机动性。采用瑞典博福斯40mm高射炮作为制式中口径高射炮 编组成预备高炮部队 可以方便地调动到最需要的地方 执行要地防空任务 充分利用现有的资源。至于师一级的野战防空 则采用20mm机关炮。历史上中国进口的20mm机关炮有瑞士厄利空、索罗通 意大利布雷达 丹麦麦德森四个类型 都是用15~20发的弹匣供弹 持续射击能力很差。应选择最新的厄利空20mm机关炮 采用60发或更大的弹鼓 提升持续射击能力。它的重量还不到300kg 完全可以由马匹驮载 跟上步兵的行进。除了防空 还能作为反坦克武器的补充 打击装甲目标。4. 大口径机枪由于财力有限 中国军队的高射炮数量不可能太多 一线步兵还需要一些更便宜 更轻便的武器来补充防空力量。大口径机枪一般都会设计成高平两用 既能对付空中目标 也能对付地面目标 而且重量也不大 是非常实用的武器。30年代典型的大口径机枪主要有美国勃朗宁M2式12.7mm机枪和法国哈奇开斯13.2mm机枪。论性能 显然是美国勃朗宁M2式要领先很多。该枪大量装备美国军队 服役了近百年也不见落后 至今还活跃在世界各个战场 丝毫没有要退役的迹象 这是最好的证明。有网友会说 30年代美国孤立主义盛行 对外实行武器禁运政策 无法采购M2大口径机枪。事实上 比利时FN公司和勃朗宁有着长期的合作关系 从30年代开始就生产M2大口径机枪。中国可以从比利时进口该机枪 完全不受当时美国的限制。因此 中国应选择勃朗宁M2式12.7mm大口径机枪 装备在团一级 不仅能作为轻型防空武器 也能作为一种反坦克武器使用。（总结）综上所述 抗战前的30年代 有两套制式武器配置方案 1. 国军制式武器优化方案如下：（有能力仿制的武器）：步枪弹：7mm毛瑟步枪弹步枪：巩造98式（或G98）（长枪管 改用7mm毛瑟步枪弹）重机枪：马克沁MG08（改用7mm毛瑟步枪弹）轻机枪：比利时勃朗宁FN D（改用7mm毛瑟步枪弹）手枪弹：9mm帕拉贝鲁姆手枪弹冲锋枪：德国伯格曼MP18手枪：勃朗宁M1935枪榴弹筒：40mm 配属步枪迫击炮：60mm 82mm 120mm山炮：博福斯M1930式75mm山炮（需要进口的武器）：野炮：德国le. FK 16式75mm野炮榴弹炮：德国le. FH 18式105mm榴弹炮反坦克炮：奥地利百禄B?hler式47mm反坦克炮反坦克枪：德国毛瑟M1918式13.2mm反坦克枪中口径高射炮：瑞典博福斯40mm高射炮小口径高射炮：瑞士厄利空20mm高射炮大口径机枪：勃朗宁M2式12.7mm机枪2. 国军制式武器备选方案如下：（有能力仿制的武器）：步枪弹：6.5mm有坂弹步枪：三八式步枪机枪弹：7.92mm毛瑟弹重机枪：马克沁MG08轻机枪：捷克ZB26冲锋枪：德国伯格曼MP18（使用7.63mm毛瑟手枪弹）战斗手枪：盒子炮（使用7.63mm毛瑟手枪弹）自卫手枪：勃朗宁M1903（使用9mm勃朗宁手枪弹）枪榴弹筒：40mm 配属步枪迫击炮：60mm 82mm 120mm山炮：博福斯M1930式75mm山炮（需要进口的武器）：野炮：德国le. FK 16式75mm野炮榴弹炮：德国le. FH 18式105mm榴弹炮反坦克炮：奥地利百禄B?hler式47mm反坦克炮反坦克枪：德国毛瑟M1918式13.2mm反坦克枪中口径高射炮：瑞典博福斯40mm高射炮小口径高射炮：瑞士厄利空20mm高射炮大口径机枪：勃朗宁M2式12.7mm机枪|http://www.360doc.com/content/15/0104/14/13530469_438086805.shtml|2015-01-04
其他媒体|1603995461|163|网易文化论坛-大陆明星|ZHO|2015-01-10 00:40:01|LOL的远程英雄大全 - 网络游戏一出戏|"神魔大陆加速器哪一款好     0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""黑暗之女安妮"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""流浪法师瑞兹"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""复仇焰魂布兰德"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""策士统领斯维因"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""光辉女郎拉克丝"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""末日使者费德提克"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""堕落天使莫甘娜"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""死亡颂唱者卡尔萨斯 "" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""冰晶凤凰艾尼维亚"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""猩红收割者弗拉基米尔"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""卡牌大师崔斯特"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""cf美服官网探险家伊泽瑞尔 "" src=""http://www.pk38.com/      0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""法外狂徒格雷福斯"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""暗夜猎手薇恩"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""皮城女警凯特琳"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""赏金猎人厄运小姐"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""麦林炮手崔丝塔娜 "" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""英勇投弹手库奇"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""未来守护者杰斯"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""狂野女猎手奈德丽"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""迅捷斥候提莫"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""寒冰射手艾希"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""爆破鬼才吉格斯"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""大发明家黑默丁格"" src=""http://www.pk38.com/      0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""琴瑟仙女娑娜"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""仙灵女巫璐璐"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""天启者卡尔玛"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""邪恶小法师维迦"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""风暴之怒迦娜"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""狂暴之心凯南"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""时光守护者基兰"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""众星之子索拉卡"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""魔蛇之拥卡西奥佩娅"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""九尾狐阿狸"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""诡术妖姬乐芙兰"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""发条魔灵奥莉安娜"" src=""http://www.pk38.com/      0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""机械先驱维克托"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""龙血武姬希瓦娜"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""远古巫灵泽拉斯"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""首领之傲厄加特"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""战争女神希维尔"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""审判天使凯尔"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""瘟疫之源图奇"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""深渊巨口克格莫"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""虚空先知玛尔扎哈"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""荆棘之兴婕拉"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""暗黑元首辛德拉"" src=""http://www.pk38.com/  0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""蜘蛛女王伊莉丝"" src=""http://www.pk38.com/      0 && image.height>0){if(image.width>=700){this.width=700;this.height=image.height*700/image.width;}}"" alt=""唤潮鲛姬娜美"" src=""http://www.pk38.com/         台服Rift玩家为你展示伊莎贝拉公主真容"|http://bbs.ent.163.com/bbs/dalustar/492561627.html|2015-01-10
其他媒体|1604667725|zhidao_baidu|生活|ZHO|2015-01-10 14:35:02|雷凌1.6自动精英好还是起亚k3 GLS AT||http://zhidao.baidu.com/question/520146340009539165.html?entry=qb_browse_default|2015-01-10
其他媒体|1604680004|meizu|综合讨论区|ZHO|2015-01-10 14:47:03|怎么煲耳机！长编煲耳机文章！|"只用港货 中级会员   一、煲机的概念及机理新耳塞、新耳机购入以后 一定很想让新耳塞和耳机发挥最大的效用来满足自己的耳朵。于是煲机成为老鸟玩家级的自然而然的选择 但是关于该煲还是不该煲的争论一直在继续。笔者借用技术和经济的角度进行简单说明。支持煲机方：新耳塞和新耳机买回来以后需要进行后期的调试和声音的再加工也就是需要进行煲机 让震膜变的松弛 从而表现出更好的声音来。反对煲机方：新耳塞和新耳机买回来以后只要保持正常的收听就可以了 完全没有必要多此一举来进行所谓的“煲”机。进行煲机的话一来没有多大的作用 二来又损伤了震膜 可谓是得不偿失。这样看来公说公有理 婆说婆有理。新手上路的话真不知道是该听谁的好 刹是迷惑。本来买了新耳塞新耳机是件愉快的事情 结果反而因为煲不煲机的问题而烦恼就大大影响了喜悦的心情。那结果是煲还是不能煲呢？假设可以煲的话新手如何操作呢？煲机有什么道理？种种疑问笔者尝试进行简单的分析和说明．笔者还是刚接触这些的时候也同样遇到了以上的问题。最开始笔者坚信新耳塞新耳机不需要进行所谓的煲机 直接正常的收听就可以了。随着笔者所见和所闻多起来 发现新耳塞新耳机还真的需要进行一定的煲机处理 这样能发挥耳塞和耳机的全部潜能 从而更加满足耳朵的需要 当然这个过程需要掌握一个度。笔者亮出自己的观点是：新耳塞和新耳机需要进行“煲”。煲好以后新耳塞和耳机各项性能逐渐稳定 指标也基本上达到了最佳 也就是所谓的煲透了。当然煲机要讲究科学不是胡乱来的。科学和谬误只在一步之间。胡乱“煲”对耳塞和耳机来说是一种极大的伤害 不仅不会发挥潜能 反而是蹂躏 由此震膜会严重受伤 直至报废。科学的煲机是磨合 新耳塞新耳机振膜折环机械顺性差 磨合经过一段时间后 顺性逐渐变好 潜能就表现出来了。这个煲机从技术角度来说恰好就是折旧 煲机怎么折旧？笔者详细说说。技术上所说的折旧其实一种设备的损耗。当然这个损耗包括有形的和无形的。煲耳塞耳机只是其中的有形损耗的层面 折旧是大概念 煲机是小概念。有形损耗又称物理损耗 设备使用是在力的作用下 各个部分受到摩擦、冲击、震动、或疲劳 最终使的设备实体受到损伤。耳塞和耳机就是“设备” 力就是电流给予震膜的作用。所以耳塞和耳机本身也是有使用寿命的。但是千万别误解了损伤 表面上看损伤都是不好的 但是有时候的损伤对设备也有利的 就是磨合过程以后就是如此。耳塞和耳机在使用中有形的损耗大致有三个阶段。图中的I期为初期损耗阶段 这一时间段很短 设备的震膜在此期间经过相对运动冲击和疲劳 很快就会把不同的发音单元进行磨去 损耗量在三个阶段中是很大的。图中的II期为正常损耗阶段 这一时期将持续很长时间 是三阶段中时间最长的时间 震膜的磨损趋于平缓 损失的部分缓慢 是震膜最佳的运动时间 基本上是随着时间做均匀的缓慢运动 这一阶段将保持状态的相对平衡 因此是比较稳定的。图中III为剧烈损耗阶段 这一阶段中 震膜的损耗度已经超过一定的限度 正常的损耗关系被破坏 此时的工作状态和情况都比较恶劣 随着时间的增加恶化的表现比较突出 损耗量是三阶段中最大的 震膜的精度、性能、幅度都大大受影响 基本上是告老还乡的时间了 基本上这一时期的耳塞和耳机已经是破音加失真甚至无法出声 已经出现了报废的表现。新耳塞新耳机进行正确煲机 就是加速其震膜“老化”的过程使的其在最短的时间内度过磨损的时期 经过“煲”的非自然力的驱使 从而提高了第二阶段的时间 使得耳塞耳机的水平提高显著并且长期保持住这个水平。特别是有的新耳塞和耳机震膜采用特殊的材料 耐冲击耐震动耐疲劳 在一段很长的时间被都不能发出好声 平常自然听可能听坏了都不能使的耳塞和耳机的能力体现出来 对于这种类型的耳塞和耳机更加应该采取煲机的处理 一旦度过这个磨合期 耳塞和耳机的表现会有质的飞跃。煲透的耳塞耳机 正常使用其性能都大大改善 而未经过煲机的耳塞耳机在自然听状态下 也有在第二阶段的某一时期出现声音的飞跃 不过这个时间是短暂而急促的 之后耳塞和耳机的素质会走下坡路。在图中分别用两条曲线来体现煲与未煲之间的区别。煲过的耳塞耳机见红色实线的曲线；未煲的耳塞耳机见蓝色虚线的曲线。二、初识白噪音白噪音、粉红噪音、褐色噪音：是由光波的谱线图就是光谱图类比而来区分这些噪音的。[白噪音]所谓白噪音是指一段声音中的频率分量的功率在整个可听范围（0～20KHZ）内都是均匀的。由于人耳对高频敏感一点这种声音听上去是很躁耳的沙沙声。白噪声是一种无规噪声 它的瞬时值是随机变化的。它的幅值对时间的分布满足正态分布。它具有连续的噪声谱 包含有各种频率成分的噪声。它的功率谱密度与频率无关 几个频率能量的分布是均匀的。它的等带宽输出的能量是相等的。它在线性坐标中 输出是一根平行与横坐标的直线。在对数坐标中 输出是按每倍频程带宽增加3dB的斜率而上升的。在人耳可听的频率范围内 具有相同能量的噪声称为白噪声。白噪声广泛用于环境声学测量中。所以从频谱仪的图形上看 白噪声在全频谱内是一条平直的线[粉红噪音]粉红噪音是自然界最常见的噪音 简单说来 粉红噪声的频率分量功率主要分布在中低频段。粉红噪声从人耳中听到的是平直的频率响应——“非常悦耳的一种噪声”最常用于进行声学测试的声音。从波形角度看 粉红噪声是分形的 在一定的范围内音频数据具有相同或类似的能量。粉红噪声的电平从低频向高频不断衰减 其幅度与频率成反比(1/f)。其幅度每倍频程(一个8度)下降3dB。噪声能量在每倍频程内是相等的。所以从频谱仪的图形上看 粉红噪声是在一个小段频谱内平直的线 并且以其倍数频率向下衰减。即1倍频 2倍频……频率越高谱线高度越低。[褐色噪音]褐色噪音的频率分量功率主要集中在低频段。其能量下降曲线为1/f^2 其波形是非常自相似的。整体来说有点跟工厂里面的“轰轰隆隆”的背景声相似。煲机就是运用收音机的白噪声和粉红噪声 根据他们的特性进行间断的煲机。新耳塞耳机初期可以采用调到无台状态下 音量偏小为宜。保持5小时以上8小时以上的连续煲机 根据耳塞耳机的不同 一般来说3天到5天时间就足够了。然后是调到有清楚的台进行第二阶段的煲机这个过程可能持续的比较长 控制在正常音量或稍大音量 有可能是一个星期或者两个星期 甚至一个月的时间。完成两阶段以后 耳塞耳机在你手里基本上已经煲的差不多了。这样操作下来 新耳塞耳机已经可以保持比较好的状态了 能尽心尽力为用户服务了三、慢煲出好声煲机的话题由来已久 众说纷纭 各有其论。老犬首次出贴怎么就来了这么个题目 实有“陈谷子烂糠”之嫌 不过“旧瓶装新酒”古今有之。诸位不妨小酌三杯 品品其中别样滋味。大凡有车族都有新车磨合的经历 何为磨合？音响行话——“煲”也。汽车的磨合可是有严格规定的 引擎要空转多少个小时 一档、二档、三档……要行走多少公里等等不一而足。为了限制新车的出力有的还安装了限速器 限制进入汽缸的燃气量 让你想快都快不了 只能在磨合完之后 才允许折除。当你磨合结束更换机油时 你才发现 好家伙！原来这油中竟有这许多残兵游勇、金属碎屑 足足吓你一个大跳。车子磨合的好坏对今后的出力和寿命的影响实在是太大了 所以凡有经验者都会延长这个磨合期限。钢筋铁骨的家伙开始竟要这般伺候 想想我们的音响器材 尤其是我们那么娇贵的耳机应该怎样去煲？煲耳机主要是煲耳机的振膜 就目前而言 静电耳机振膜的厚度已薄到1•35微米 动圈耳机的振膜也只有几微米到十几微米（我们头发的直径大约是60～90微米）。振膜本身在制造过程中就存在内部应力 在粘结音圈和固定在骨架上时又产生了装配应力 我们所说的煲耳机就是使这些应力逐步消失 使振膜逐步顺化发出好声的过程。我常看到一些Hi-Fi大师们的器材试听报告 水平高低且不评论 只是那开头大多是先把器材开足马力猛煲它三天三夜 让它受尽皮肉之苦 自以为进入佳境 而后才是如何如何好声好声评论一番。天长日久煲机之法由此而生 效仿者不计其数。如此煲法就不怕损伤器材 落下隐患 好声不长！我以为音响器材虽不是工程机械、铁车钢马 但也有相通之处。好事需多磨 慢煲出好声！煲机还是分为舒筋、通络、习武、打擂、出道五步为好。以耳机为例：1、舒筋——使用正常听音强度三分之一的音量驱动耳机12小时（用100～1500Hz/5s扫频信号更好）；2、通络——使用正常听音强度三分之二的音量驱动耳机12小时（用50～1800Hz/3s扫频信号更好）；3、习武——使用正常听音强度驱动耳机72小时（用20～20000Hz/2s扫频信号更好）；4、打擂——使用正常听音强度三分之四的音量驱动耳机24小时（用18～2200Hz/1s扫频信号更好）；5、 出道——进入正常使用阶段。我想这种煲机方法最少有两大好处 第一可以了解煲机各阶段音质变化的规律 理解煲机的作用 积累经验；第二可提高器材性能 不留隐患延长器材寿命四、怎么煲耳机 让声音听起来更美妙！随身听爱好者们常常会拥有一副好的耳塞 但在开始使用时发现并没有像其他人谈论的这么好 难道是自己买到了假货？非也！其实那是因为没有进行购买后的第一道工序——“煲”。为什么要“煲”耳塞其实在音响界 很多东西都需要“煲”。包括音源、功放、音箱等等。所谓的“煲”就是让这些东西运作一段时间 以达到最佳的效果。我们刚买回来的耳塞 不出意外的话都应该是刚出厂的产品。这些耳塞从生产线上下来的时候 震膜一次都没有用过 因而会很硬。这种情况下的震膜突然震动起来 会感觉很不自在 声音也会略微走样。如果一开始就好好的“煲”一下耳塞 那么就会把它的震膜逐渐弄松 这样再听音乐时 震膜震动起来就会非常的自如 音质也较先前提高不少。“煲”耳塞前的准备其实“煲”耳塞（机）并不困难 但是需要时间和一定的技巧。首先 你需要一个可用来长时间放音的音源。因为“煲”耳塞可不是一会儿半会儿的事情 有时候甚至需要100个小时以上。其次音源中要有频响范围很宽、动态效果舒缓、层次清晰、高中低音各成分适中的音乐有这样效果的音乐要比一般音乐“煲”起来效果更明显。还有一点就是音源输出功率一定要够大 而且要和用户的耳塞档次匹配。比如要“煲”HD580就不能用普通随身听 随身听可能连推都推不动 还怎么让震膜松动呢？一般来说 随身听只适合耳塞和一些低阻抗耳机使用。一般而言 如用电脑声卡和收音机“煲”耳塞的话 需要比较长一点的时间。而用输出功率很大的CD随身听来“煲” 时间要短一些。“煲”耳塞的操作首先 我们需要数张CD碟 这是因为CD音质是目前民用级别（撇开并不实用的SACD和DVD-AUDIO）可以达到最好效果的音乐质量 而且碟片相对来说比较便宜 以下所有操作也均以CD随身听为例。“煲”机碟最好是张频响范围非常宽广的碟片 单独使用一般的纯人声碟肯定不行。推荐一些正版的发烧碟 比如《TITANIC》、《阿姐鼓》和《1812序曲》等等。还有一些优秀的流行音乐和中国民乐也是很不错的选择。下面笔者就来“煲”好你的耳塞。《TITANIC》电影原声CD中的第3段《SOUNTHAMPTON》、第9段《THE SINKING》和第10段《DEATH OF TITANIC》。《SOUTHAMPTON》虽有抄袭贝多芬的《欢乐颂》之嫌 但声音层次非常分明 乐曲包含的信息量也很丰富。高中音柔顺致密 隐隐而来的阵阵低频能量予人一种深邃感。这首曲目在全频段都有突出表现 对于耳塞的全面震动是非常有好处的。而《THE SINKING》和《DEATH OF TITANIC》除了与上面一首有同样出色的全频表现以外 在动态上更胜一筹 整体声音能量十足 如果没有“煲”就听这样的曲子 耳塞的震膜要“受苦”了！国产动画电影《宝莲灯》电影原声CD中的第4段《序曲：宝莲灯》和第13段《望月节的舞蹈》。《序曲：宝莲灯》一开始声音较为轻柔 但越到后来 声音动态越大 能量也越多。中间还夹杂着一些人声的合唱 应该说是非常不错的曲子 唯独其低音略微少了一些。《望月节的舞曲》中一开声的低频以及中间一段女声对于耳塞中低频的提高都很有帮助。《滚石24K24BIT金碟--万芳》CD中的第一段《猜心》是笔者用作试音的保留曲目 用来“煲”耳塞也是非常不错的选择。这首曲目的第一段主要是人声独唱 不过到了后面 乐器就越来越丰富 但整体仍可算是轻柔。“煲”耳塞不能一直用大动态来“煲” 也需要在中间做一些调整。而且 这首曲目中的人声非常出色 可以用作“煲”耳塞结束以后的试听之用。其实优秀的曲目太多了 笔者在这里推荐的只不过是冰山一角而已！把随身听和耳塞准备好 放入碟片 音量上要开的大一些。现在的随身听为了延长播放的时间 输出功率普遍较低 用户大可以把音量开到90%以上 不过最好不要开效果！“煲”耳塞的过程中要一步一步的来 首先用一些舒缓的音乐 比如上问中提到的《猜心》 先放5－10个小时。然后再换略微""厉害""一点的音乐 如《SOUTHAMPTON》 继续播放10小时以上 最后才是诸如《THE SINKING》和《DEATHOF TITANIC》之类的音乐 一直要播放到耳塞基本上“煲”好。为了确定耳塞“煲”的情况 用户可以每隔10小时听一次 一般来说 效果都会有一些差距 等到差距不明显的时候 就可算是“煲”好了。当然 这种鉴别方法也不是很容易实现 那么就准备“煲”50~100个小时好了。不过要达到大功告成就需要日常不断的使用才行 要使耳塞真正达到最佳效果 时间上一般需要2个月左右。前后声音的对比：笔者“煲”耳塞“煲”过很多 最有感触的就是索尼（SONY）MDR-E888了。这是一款目前相当高级的耳机 市售价在人民币400元左右。但是这款耳塞刚买回来试听的时候 常常都会有高音发干 中频毛刺多多等问题 让人觉得完全不值400大元。不过一旦MDR-E888“煲”好了 那么她就会放射出耀眼的光芒：柔顺的高频、温暖但绝无毛刺的中频、深沉有力的低频 简直不敢相信是同一个耳塞。个人认为 MDR-E888是笔者见过的耳塞中最需要“煲”的一款 这可能和它独特的生物震膜有关系。其它的耳塞也都需要“煲” “煲”过以后都主要体现在低频弹性感得到加强 高频柔顺感有了提高 只是结果好象没有MDR-E888那么夸张！“煲”耳塞是一个漫长的过程 需要将“煲”和日常合理使用相结合 如果能正确的“煲”好你的耳塞 那么 相信她一定会给你带来不一样的惊喜！五、测试&欣赏天碟荟萃前言：市面上的音箱、耳机品牌繁多 让人眼花缭乱。简单地看一些评测、推荐不失为一种省心、省力的作法 但真正要选购到您心仪的、适合自己口味的产品 还是坚持“耳朵收货”的原则为上！本文将介绍几张有口皆碑的天碟 它们不但适用于测试、选购 也是音乐欣赏的上上之选；同时考虑到电脑玩家的口味、多媒体电声产品性能的局限性等因素并没有推荐那些较难理解的古典天碟。需要注意的是 由于个人喜好、水平等限制 这些CD也最多只能算是音乐天堂中的沧海一粟而已 正所谓没有一张榜单能尽收天下铭器 本文也难免挂一漏万 希望大家理解。中频人声：有句发烧俗语曰：“人声是肉。” 对于价格便宜的设备来说中频是否耐听显得尤其重要（追求高低频的延伸与质感、解析度并不现实）。同时 人声也被称作最难表现的乐器 所以本次推荐以人声为主。女声：1.蔡琴《机遇-淡水小镇》蔡姐相信已没有多作介绍的必要 其老歌是发烧友、爱乐者人手一张的必备之物。该碟的钢琴伴奏和编曲皆由音乐奇才鲍比达一手包办 洋溢着让人如痴如醉的诗情画意。正如该专辑的名字一般 《机遇》自始至终带给人的却是一种真正的音乐享受 让人轻易进入那散发着淡淡幽香的音乐隧道……当然从纯Hi-Fi角度看《机遇》也是一张不可多得天碟 无论是蔡姐的浅吟低唱还是鲍比达一手清新脱俗的钢琴都无可挑剔 人声的质感、口型 钢琴的巨大共鸣、弹跳感 静谧的背景和深广的音场等等 皆为上成。推荐：Track1“机遇”（考验人声）、Track6“月光小夜曲”（考验人声及音频系统的透明度、纯净度 音场的深度、广度）等。记得《机遇》在第六届国产音响展上几乎被放“滥”了 原因没有别的 只因为它把音乐和音响这两个因素结合的是那么完美。2.朱哲琴《阿姐鼓》《阿姐鼓》是由何训田作曲 何训友作词 朱哲琴演唱 上海音像公司于1995年出版 是国产CD中不可多得发烧天碟。作者曾历时二年多 亲赴** 走访寺庙 深入藏民基层 在仔细观察雪山、草地后完成了这部发自内心深处的巨作《阿姐鼓》。该专辑共由7首曲子组成 制造精良 纤细处丝丝入扣尽显女性的柔美 高亢处宏伟壮丽如同**一望无际的蓝天。朱哲琴的嗓音婉转飘逸 “没有阴影的家园 没有阴影的树 ……”歌声仿佛已将我们带到世界屋脊那纯净、神秘的世界！该碟不但人声极其出色 低频也是雄浑厚实下潜很深 就像世界屋脊的高海拔带来的压抑感觉一样。《阿姐鼓》并非浪得虚名 不信您大可跑到音响店瞧瞧 也许试机时店员就会放进一张《阿姐鼓》以“炫耀”低频哦！优秀的女声天碟还有许多 像王菲《天空》、Loreena McKennitt《神迷之书》、杨小琳《禧乐》、戴安娜.克劳《When I Look In your eyes》、沙拉.布莱曼《月亮女神》等等。男声：1.腾格尔《天堂》蒙古族歌手滕格尔有着大漠男儿的豪迈和热情 他的人声中气十足、爆发力极强 也是音响店试机的常用CD之一 一般中高频不过硬的系统被腾格尔一嗓子就会吼的洋相百出。这次推荐的是其XRCD2版 音效较《四十独白》大有提升 中国联合交响乐团的伴奏也增添了更多细节和更雄伟的场面。这是近年国内乐坛不可多得的精品音乐集 歌唱者的沧桑、成熟、热情值得品味。2.《阿淘的歌》阿淘本名陈永淘 是台湾新竹的一位客家民歌手。无论是歌唱者还是出版商都可谓默默无闻 但《阿淘的歌》何以被专业媒体冠为“近年少见的男声试音典范”呢？！有两个原因 一是感人至深的演唱。15首歌曲全部由阿淘自己作词作曲 他的演唱很真诚 很自然 毫无修饰做作 嗓音中流露出一种沧桑感但却又不乏积极向上的因素 与《机遇》相似 《阿淘的歌》也是以平淡感人取胜 这也许正应了“平平淡淡才是真”这句老话吧。其次 该碟的录音漂亮到无懈可击 看看《音响世界》是怎么评价的吧：“《阿淘的歌》录音非常漂亮 绝对是近年来男声发烧录音的典范 假如在大型视听欣赏会中采用 相信它一定会有镇场的效果……最适合校验Hi-Fi组合的音场还原能力……”相信听完本碟 会激起您对音乐、生活的无限热爱 如果只用来试音确实就太浪费了。推荐：《仰葛煞》、《春水》、《想问》、《日出部落》等。3.中国八只眼《青叶城之恋》也许本碟在录音和包装方面比其它几张CD没什么优势甚至稍差 但是真正重要的是它会带给您前所未有的舒适音乐感受。八只眼男声四重唱演唱形式轻松、活泼 演唱曲目兼顾中外民歌风采 在声音运用上把传统、民族和通俗唱法融为一炉 使一首首名曲老歌丰满深沉、欢愉浪漫 散发出极强的艺术魅力。同时录音水平在国内也算优秀之作 整体定位清晰、层次较好、空间感出色。《三百六十五里路》、《弹起我心爱的土琵琶》、《同一首歌》、《游击队歌》、《大坂城的姑娘》等等大家熟悉的经典歌曲获得重生 是一张雅俗共赏的优秀CD。此外值得购买的还有意大利瞎子男高音Andrea Bocelli的最新大碟《CIELI DI TOSCANA》、夏韶声《谙》、飞鹰乐队《加州旅馆》、世界三大男高音作品等等。高频：1.吕思清《四季》维瓦尔第的《四季》号称再版次数最多的古典名曲 我国小提琴顶级大师吕思清用6把价值上亿的名琴再次演绎并由马可波罗公司以顶级录音器材精心打造。在世界乐坛享有盛誉的中国小提琴家吕思清加上The Stradivari Society（斯特拉迪瓦里收藏协会）提供的6把绝世名琴 并由世界一流器材、录音师录下这辑发烧级“四季” 是发烧乐迷绝对值得收藏的天碟。听完此碟 如果您的音频系统足够强劲相信就会大致明白成天挂在发烧友嘴边的“天碟”是何含义了：无论是高频区的解析力、延伸度还是乐队整体的定位、层次都堪称示范级水准！不过由于该碟解析力极高、透明度非常好 所以能把它放过关的普通设备可谓寥寥无几了。推荐试听片段：春（第一乐章）不建议选择吕思清的《四季》）2. 阿卡多《Diabolus IN Musica》（魔鬼小提琴）该碟由意大利著名小提琴家阿卡多演绎 帕克尼尼的经典作品收录了不少。在音响店这也是一张“不敢”随意乱试的天碟 普通低价器材放出来的声音索然无味 全无感觉……Track2《La Campanella》也叫“Ensemble”（帝王） 由阿卡多拉来犹如天外来音一般 小提琴的松香味、木质感、擦弦等等如实奉上 余音绕梁三日而不绝！好的音频系统重放本碟让你根本感觉不到音箱的存在 而在两个音箱中间则可以“看”到一把名琴在飞舞……对自己的听音设备很满意的朋友不妨试试本碟 也许您会有新的认识。推荐：Track2《La Campanella》、Track3《Capriccio per violino solo n.5》低频／整体：由于成本的限制 多媒体音箱的低频不可能有什么“力水” 而同价位的耳机则要在这方面好上不少；加上低音单元的尺寸限制 个人认为在多媒体音箱上低频的质远比量重要的多！而中低价位耳机缺乏的则是真正的低频下潜 厂商一般会人为提升低频作为“补偿” 使他们的产品听起来也有那么点“震撼人心”的意思。3.Telarc唱片公司《1812序曲》（DSD技术录音新版）可以肯定的是目前市场能将《1812序曲》摆平的Hi-Fi系统非常少 但考虑到它的“权威性”还是做一推荐。1812序曲是俄罗斯著名作曲家Tchaikovsky（柴科夫斯基）最出名的交响乐作品之一 录有真实的炮声 足有摧毁器材的魄力！因此大家播放此碟前一定要设置安全的音量 免得“机毁人亡”！康泽尔指挥下的辛辛那提通俗乐团演奏老练出色 音乐感强烈。新版本的《1812》不但管弦乐部分极其出彩而且人声合唱部分一流 是一张不可多得的试机天碟 也难怪那么多的器材发烧友将其作为“看家”之作了！4.阎学敏《炎黄第一鼓》也是音响界试音的必备软件之一 荟萃了中国鼓韵文化的精粹 以巧妙的手法展现出一幅华夏人民的生活风貌。《鼓诗》在国内音响界早已是公认的低频天碟 系统的低频到底如何 一试便知！如果试听时感觉低频力度好、速度正确、鼓皮的涨力都仿佛历历在目 同时也没有什么发散、发蒙的感觉 那么系统的低频基本就过关了；如果能“看”到鼓皮的颤动、阎学敏手起棍落的爽朗那么真该羡慕您才对……5.雨果《雨果发烧碟8》这是一张很常见的发烧碟 采用24K金压片技术 加上HDCD技术的辅佐 使得该碟音质不俗。Track1《大黄河》动态惊人 气势极大 用来考验音箱的动态再好不过；Track2《在那遥远的地方》为杨小琳的个人“show” 她那迷人的嗓音以及悠远开扬的风格让人百听不厌；Track9《阳春白雪》有着近似打击乐的奇特效果 同时爆棚场面也是耐人寻味……总之 这是一张适合发烧友及民乐爱好者的大碟 不容错过。6.《拿索斯发烧「骚」》最后出场的是来自以性价比高而著称的拿索斯 是该公司在过往十五年来所灌录的发烧录音的一次大汇演。此碟所辑录的曲目皆是权威音响杂志主编的精心推介 其中包括国际权威音响天书美国杂志《绝对音响》（The Absolute Sound）、誉满大中华地区的两本权威音响杂志《音响技术》（Audiotechnique）及《发烧音响》（Audiophile）与响誉全球的音乐音响英国杂志《留声机》（Gramophone）。《拿索斯发烧「骚」》网罗音响示范级佳作 古典音乐精华尽收本碟。交响乐气势恢宏无比 录音效果令人瞠目。六、避免低级错误:褒耳机的种种致命做法注意：这里讨论的耳机范围不包括顶级发烧级别 只是给初步入门用户的参考。如今 越来越多的人已经了解到耳机对于音质改善的重要作用 无论是接随身听还是声卡 许多人都在研究升级购买高档耳机来体验“HI-FI感觉” 要知道 欧美真正的有钱人都是玩音响的 几十万的大家伙买不起至少要弄个好耳机来享受享受吧！但越是高档的新耳机越要细心褒 因为震膜在这个时候还没有舒张开 紧绷绷的 出来的声音也很令人失望 一般的表现是高音刺耳 中频干涩 低频缺乏细节 要经过一段时间（大约200-400小时）的放音、也就是“褒机”之后才能“逐渐”体会到革命性的变化（注意 是“逐渐” 这个过程很激动人心的 就像《角斗士》电影里的拉塞尔•克劳越来越强壮的性格和身体） 相关的介绍在网站和平面媒体上都已经很多 这里要重点说的是一些常见而致命的错误。在跟一个资深音响人士聊天时他说 现在返修的很多耳机都是在褒机的时候方法不当坏掉的 “要是方法得当 褒好以后正常情况下几年也不会坏的。” 又说到一个很夸张的例子 一个自称是“清华大学”的用户买了一个几百元的耳机回去以后 用电脑上的“频率发生器”产生20Hz的声音 然后用耳机接声卡试听 要“褒低频” 并且看看耳机究竟能不能达到标称的20Hz下限值！当然结果是耳机拿回来修了。他们特意就此写了警示文章 摘引：“在这里我们想请读者注意 20Hz是人类的听音极限 就是说在20Hz时人类的耳朵刚刚开始有知觉（肯定还有一部分人根本就听不到） 在20Hz的情况下人耳朵的灵敏度极低 要使耳朵听到声音 势必要使之振幅极大。在这种情况下 小小的的耳机怎么能不打底 又怎么能承受得了。因此读者应记住千万不要用这种方法来试验耳机 这是十分错误和有害的。举例来说人耳对3000Hz的灵敏度与对20Hz时的灵敏度会相差20～80dB|我们知道灵敏度每相差3dB推动功率就差两倍 同样的 差6dB就差4倍 差9dB就差8倍。那读者估算一下如果你要听到20Hz要输入多大的功率？而且20Hz的信号势必要使震膜的振幅极大、同时音圈的阻抗降低 电流急剧升高 使音圈发热变形 进一步导致震膜变形 造成破声、蹭圈等永久性破坏 即使是短时间的试听也会使音圈打底的。”同样 用一些频率发生软件来褒耳机也是很危险的 固定频率的强电流轰击很容易损坏新耳机舒张度不够的震膜。前阵有个网友在QQ上求救 说他的一个400元的耳塞出现破音了 我说你是不是用软件褒来着 他说对啊你怎么知道啊 我都褒了2个多小时了……。——如果说这些专业的软件有用的话 那只能是专业音响技术员用适当的方法很小心地在特定的设置、输出功率和时间等等因素综合下 对耳机的“磨练” 普通用户如果用这种工具 一不小心就会弄坏耳机 即使是使用了很久的旧设备在这样的“折磨”下也可能挂掉 更不要说脆弱的新耳机了！此外 也有许多人喜欢用强劲的音乐来褒 比如重金属摇滚、电子舞曲 而且开很大音量 这同样会很快造成耳机夭折或产生噪音。特别是如果刚打开包装便用大音量强音轰击 那么即使是素质很好的耳机单元也受不了。——只有在完全褒开以后 能够承受的“磨砺”就相当大了。唯一普遍适用的褒耳机方法是“渐进” 刚开始用轻柔一些的音乐 在较低音量下让耳机先舒缓10-30小时 然后用普通的音乐（摇滚、舞曲除外）在中等音量状态褒100-200小时；如果这时你听着高音不刺耳了 变得圆润自然 中音温暖亲切 低频再也不是混成一团的轰隆隆 而充满细节 那就恭喜 OK了 绝对不能急功近利。"|http://bbs.meizu.cn/thread-5466805-1-1.html|2015-01-10
其他电视|1617181564|cztv|zhejiang|ZHO|2015-01-18 22:11:01|杭州赏腊梅正当时 2015杭州赏梅全攻略|2015-01-18 09:07 来源：杭州网  -->  　　孤山的蜡梅 记者 许康平 摄昨天上午 一则“2015杭州赏梅全攻略”在网上热传。又逢杭城赏梅时 眼下的梅花开得怎么样了？昨天 快报记者先去植物园和孤山看了看。“要看梅花还早嘞 都还是些小花骨朵呢。进去看看蜡梅吧 黄颜色的 开得正旺 味道也清香！”下午 刚走进杭州植物园南门 就看到一位大伯笑呵呵地给几个小年轻指路。“蜡梅不就是梅花吗？”一位姑娘一脸迷茫。“当然不一样啦！”大伯对着姑娘的手机屏幕一指 “你们对着这个网上的攻略来看梅花 那可能要失望了。照片上这些红梅白梅 还没怎么开呢！”旁边一位拿着单反相机的帅哥走过来“科普”：“蜡梅是黄色的 植物学上有个单独的蜡梅科。你们想看的梅花啊 属于蔷薇科 有白的、粉的、红的 还有绿的 要看满树梅花绽放 得等春天啦！”植物园的保安朱师傅说 这几天的游客不算多 大部分是来赏梅的 而分不清楚蜡梅和梅花的 的确有不少。不过朱师傅觉得 分不清也不要紧 总归都是美丽的花 进园看看总不会失望。杭州植物园高级工程师胡中也赞同：“灵峰有1000多株蜡梅 最近一段时间竞相争艳 正是观赏的好时机。而梅花 现在虽然开得不多 但偶有几朵绽放的意境 也是很美的。所谓‘寻梅’、‘探梅’ 就是要你顺着淡淡的花香去寻寻觅觅 这才有乐趣嘛！”的确 昨天灵峰的蜡梅园和品梅苑内 清雅的花香随着寒风阵阵浮动。一株株蜡梅花开满树 凑上前细看 明黄色的花朵仿佛金雕玉镂一般 有些还裹着丝丝紫红色的花蕊 显得分外澄澈晶莹。和蜡梅相邻的一排排梅花树中 也已有几株江梅、粉红朱砂以及龙游梅有零星花朵绽放 很是可爱。对于花了不少时间才“寻”到它们的游客来说 无疑是一份惊喜 大家纷纷欢快地上前拍照。“四面有山皆入画 一年无日不看花。”对于爱赏花的杭州人来说 冬天怎么能错过赏梅呢？最近几天都是多云到晴的天气 大家不妨去西湖边走走 去植物园逛逛吧。如果你想伴着一汪湖水赏蜡梅 孤山脚下也是个不错的选择。在中山公园入口处 以及孤山公园林社旁 也有不少蜡梅吐露暗香。现在已经到了梅花争相竞开的时候 杭州周边更是有不少值得一去的赏梅胜地。我们特地为大家盘点2015年杭州周边的赏梅地！　　孤山：以梅为妻、鹤为子孤山自古便有杭州“赏梅三大胜地之首”之誉 深受杭州市民和游人的喜爱。孤山梅花始盛于中唐 有梅株遗传至宋初。南宋孤山皇家园林植梅盛极一时 凉堂、西村植梅都有数百株。孤山梅花早在唐朝就已著名 白居易在他的一首诗中就有“三年闲闷在余杭 曾为梅花醉几场 伍相庙边繁似雪 孤山园里丽如妆”等句。　　如何前往乘27路、118路、k27路、k850路、y1路、y2路、y3路、假日4旅游专线、游10线/y10到岳庙站下车 步行前往或乘西湖游船到中山公园上岸。　　灵峰：暗香浮动灵峰探梅“灵峰探梅” 位于杭州植物园内的青芝坞。五代吴越国时此地建有建有灵峰禅寺 因北宋诗人苏东坡的喜爱和题咏而出名。它和西湖孤山、西溪并称为杭州的三大赏梅胜地。1988年春 园林部门重新辟梅园四百多亩。植梅五千余株 其中有罕见的“夏腊”二百株。如今在这青山环抱 树木葱郁的幽谷中 草地如茵 梅林似海 楼阁参差 暗香浮动 景色十分诱人。　　如何前往乘15路、27路、28路、82路、807路假日旅游专线、k15路、k27路、k28路、k807路、k82路、y1路、y4路、y6路、游3路空调到玉泉站下车 步行前往。　　超山：十余里遥天映白超山的梅花以观赏“古、广、奇”三绝的梅花而著名。每当初春二月 花蕾爆发 白花平铺散玉 十余里遥天映白 如飞雪漫空 天花乱出 故有“十里香雪海”之美誉 为江南三大探梅胜地之一。中国有五大古梅。晋 隋 唐 宋 元五大古梅 超山就有其二——唐梅和宋梅。别的地方的梅花只有五瓣 惟独超山梅花却有六瓣 甚是奇怪。　　如何前往乘坐319路、786区间在超山站下车 步行前往。　　西溪：舟从梅树下 踏雪赏梅花西溪探梅在杭州西湖旅游史上也曾有过篇章 清代的“钱塘十八景” 其中就有西溪探梅。西溪主要栽植的是“绿萼梅” 明清时被称为西溪梅 是梅中极品。每到暮冬初春之时 游客便会从四面八方赶来“除旧迎新 品茗赏梅”了。“西溪探梅”最大的特点是可以摇舟作岸上观 梅树野趣天成 乘船过秋雪庵、西溪梅墅、香雪屋等处 两岸梅竹绕村 红梅白梅如云如梦 还有芦苇重重、渔翁撒网、船娘唱晚、一派田园风光……　　如何前往乘坐：193路、310路、356路、506路、k310路、y13路在周家村(西溪湿地)站下车。  返回|http://n.cztv.com/zhejiang/652079.html|2015-01-18
其他媒体|1625947205|youku|科技|ZHO|2015-01-24 01:03:01|daya550 p2飞控夜间炫彩LED悬停2|视频: daya550 p2飞控夜间炫彩LED悬停2|http://v.youku.com/v_show/id_XODc3NTk3NDY4.html|2015-01-24
기타|1626281958|newsworthknowingcn|Main RSS|ZHO|2015-01-24 09:18:01|2015-01-22|"（周四 81起）冲突＊［强征］2015.1.22 重庆市 江津区 珞璜镇用户vk33gug3i1重庆江津市珞璜政府因征地 不付农民赔尝款强行施工把七十几岁的老太婆打倒在地 这就是政府罢工 罢市＊［工人］2015.1.22 山东 德州市 德棉股份有限公司 （德州国棉厂）妙明本性#几个月不发工资出现场景#李志卫 德州市国棉一厂拖欠工人工资半年 养老保险5年不交。工人上市里讨薪 警察镇压手无寸铁老百姓 怎么不抓贪污工人工资的人。一天里也没有一名电视台记者出现 无一市政府领导说话。被逼无奈 走极端！刘莹: 浩浩荡荡几千人日谷番冬狮郎 听说国棉厂闹事了 该 我这个好奇心啊 下班路上看到火车站黑压压的一片人 各种好奇 听人家说国棉的闹事了 我去了 想拍照留念诺基亚神器不行……用户**********德州市国棉厂发生了工人游行罢工事件 O微博视频反动派 德州迎宾路德棉集团职工索要欠薪上街了|德棉一厂2000多人欠薪已4个月。到处都是井叉井车 这也是党国一贯的对待罢工工人的原则。用优势的暴力武器对待手无寸铁的工人 用最恐怖的威胁迫使工人屈服。德棉集团是德州最大棉纺公司 上市企业 拖欠社保已5年 人均1千元多点的月工资巳拖欠4一9个月。与厂方和政府多次交涉无果 忍无可忍的工友们今天走上了街头。工友们加油！（18:15）德棉一厂欠薪 工人罢工封路进行中。（18:21）目前罢工工人人数略有增加。（18:26）井叉仍是严防死守 可以走但绝不让进（18:37）最新消息 下午抓了6个人 现在已放回2人 工友鼓掌欢迎罢工已于晚7点多钟结束 历时5个小时 当局承诺先付两月工资。唉！就是这么容易糊弄。口头协议已达成 1、月底前支付两月工资 2、放了被抓的工友。现场等待放人中 党国最拿手的秋后算帐也进行中了。历时5小时轰轰烈烈开始的占路罢工就这样乱轰轰的散了。只用了5分钟的散场出卖了自己也出卖了工友的努力。也须 下午有人被抓的时候 就都盼着有人喊：“都散了吧”！这样一群心怀各异的人凑在一起还能要求什么呢！唉！！齐鲁高俊飞德棉股份有限公司员工闹罢工！！我的名字就是萌萌哒在德州也能见着游行……国棉厂不发工资……特警已把通往火车站的道路封了 现在正堵在这个路口 郭晓健_要向前这年头。国企破产 没钱发工资了 员工示威游行 连特警都出动了 年根儿了 要钱买年货啊 铠钾回趟家而已 路遇国棉厂工人罢工 人真的太多了 各种警车封锁道路啊啪啦啪啦噼里啪啦Hsss这是咋了痞子万人迷cc中国特色… 呦吼小博山东省德州市国棉厂三个月不发工资 正在闹事！ 皆有可能strive：被抓了几个YG刘运果德州人民真伟大！国棉厂工人大罢工！上海画廊-王先森德州弊端可以追溯到贪官黄胜时期.政府不作为.经济凋敝.从记事的时期起很多单位都破产工人下岗.直到现在工人无薪可拿.他们是最底层普通工人维护自己权益却被各种警围堵.某人你在不管事只吃官饭离处分也不远了天天学习好100分欠工人工资 逼的工人走这条路 小半年沒有工资了 还有好多双职工可咋活 动静大了 制止 说服 规劝。事情过后 依然是沒有结果。大TTgo （出）出事了 麦多响叮咚 在迎宾市场那里 国棉厂的罢工了lengmo_love  （19:15）就是因为这群人 他们在火车站闹 搞的我们现在还不下班 在市政府守着！fuck！你们倒是赶紧他妈的冲过来哎！全部抓走了一了白了 我们也好撤退了！shit！枯叶蝶 山东省德州市国棉厂闹事了4个月没有发工资了没有人性＊［工人］2015.1.22 广东 深圳市 宝安区 裕达富电子有限公司889开心今天差不多全厂人罢工啦 还我薪水、还我工事、加薪水咯！俊酷未来 （沙井）沙井和二裕达富电子 员工罢工。乱扣工资 辞工又不批 已经两天啦 110来了似乎也没用。罢工程序升级 在车间打架斗殴。小海马go: 今天我亲眼目睹一切 公司领导喊治安仔进来打员工 他妈的这些人简直就是畜生俺是耕田的5533 （罢工）罢工正在进行中。深圳市宝安区沙井镇河一裕达富有限责任公司 罢工还在进行中 全体员工停工放假 时间不限。有图。 侵犯农民工劳动权力 工厂血肉 有目共睹。工厂谎声按劳动法 进到工厂里 工资加班六打折 根本没有一点劳动法的规定 工厂制度只有罚没有奖。＊［客运车］2015.1.22 河南省 郑州市 巩义市Another_King两家客运公司的争执：一家要求涨价 另一家没涨 便在国道上堵路～～巩义旅游公交。 半つ人间 （这）这康百万到雪花洞的车都咋了 都被人挡这儿不让走了！你觉得你能了 刚从那路过 据说是和往米河类车路线重了 让他们换条路线 不愿意。所以就堵路了！小黑狗ac 好想不是路线重的问题 是米河类车自身的问题导致罢工 然后他们堵着雪花洞的车也不让走 不然他们的罢工就起不到作用了西皮流水830625 米河车罢工了。昨天就没有米河车跑。光有到雪花洞的车 今天就堵人家车 米河车太不像话了。罢工原因可能说是取消油补了 要求票价提高。＊［客运车］2015.1.22 黑龙江省 佳木斯市 抚远县点艹个种不服 （县）县政府被堵了！谁知道啥情况？有话说也不能让客车停运啊？百姓出行怎么办啊？跑黑车的得注意了 消停回家呆着吧 运管要抓了 抓到就得三万。喔叼腻捞姆 小客车维权 黑车确实猖狂 有些黑车主竟然狂言要干没小客车 然后他们就涨价跑＊［商户］2015.1.22 广东 广州市 荔湾区 永盛市场姚記厨神市场升租、永盛市场再一次蔬菜区罢工！俩边空空的 示威＊［工人］2015.1.22 四川 资阳市 安岳县 成安渝高速风潇水寒笑天成安渝高速公路的农民工干了活拿不到自己的血汗钱 公理何在啊…＊［工人］2015.1.22 湖南 永州市 零陵区政府玻璃窗里的苍蝇”创卫”工程款拖欠 民工集聚区政府＊［工人］2015.1.22 陕西 西安市 灞桥区 浙江驰成建设公司0MoMaek0何时归还我们血汗钱＊［工人］2015.1.22 山东电力建设第二工程公司（赞比亚项目）GXYbaby*******怒讨血汗钱 异国他乡 黑心山东电建二公司一手遮天 工资不发放 工人兄弟没吃没喝 有血性的朋友们转起来。让全世界人都看看山东电建驻赞比亚项目对工人兄弟所下的黑手＊［工人］2015.1.22 云南路桥三公司用户ie3a8kxaql云南路桥三公司农民工要不到工资 还要打人＊［工人］2015.1.22 湖北 荆州市近在咫尺的海角天涯火车站这边听说有农民工讨薪＊［工人］2015.1.22 北京市 朝阳区 金星园戴政旭Damon金星园小区门口发生一起讨薪事件 具体原因不明 大家随意感受下！＊［工人］2015.1.22 浙江 金华市我是一朵蘑菇妹纸有困难 找政府 这没错！要不到工资 找政府帮忙 这也没错！可是你总要给点时间 说点诉求 派几个代表吧！堵车 堵门口 堵公路 这也是够了！本来觉得是同情 现在却觉得真是不讲理啊！还好警察叔叔是万能的！把他们劝走了＊［工人］2015.1.22 江西 九江市 都昌县 盛世西湖（网页链接）《都昌盛世西湖楼盘农民工在县政府门口拉条幅讨薪》1月22日下午 都昌盛世西湖楼盘农民工在县政府门口拉条幅讨薪 22号上午农民工在盛世西湖工地现场讨要说法无结果后 部分农民工下午来到县政府门口拉起条幅 意欲引起相关部门的重视。条幅上声称 都昌盛世西湖拖欠民工工资2年 血汗工钱至今未还。据了解 都昌盛世西湖楼盘原开发地址的老造船厂一带 规划初期是几十亩大型社区楼盘开发 后因合伙人及其他原因拆分成多个楼盘开发 也就有了现在的盛世西湖、胜发国际等楼盘。＊［工人］2015.1.22 重庆市 巴南区baby_U_know路遇建筑工人追讨工资！人手两个饭盆儿a丫头小妮儿：我去取车时还没散 黑多警察来了在那儿 车取出来看到讨薪的人和警察都没了。怎么回事？？＊［工人］2015.1.22 黑龙江 齐齐哈尔市 广厦集团清远幽香01今天上午齐齐哈尔市政府机关大楼门前 在寒风中等待答复的讨薪农民工＊［工人］2015.1.22 浙江 杭州市 钱江开发区 钱江国际广场喻小森据说拖欠农民工工资 公安都来了。钱江开发区管委会那 钱江国际广场。＊［工人］2015.1.22 四川省 成都市 温江区开满虞美人的山坡上班途中遇见维权的他们 虽然只有下车走路到办公室 但希望他们维权成功 拿到血汗钱 回家过个开心年！ ＊［工人］2015.1.22 河北 邢台市 锦江花园漂泊人生万岁邢台市开发区锦江花园工地民工讨薪。邢台市政府门口农民讨薪现场政府部门的监管不得力 才导至农民工讨薪困难 民工真没有人权了吗？＊［工人］2015.1.22 河南 许昌县 苏桥镇 龙成集团许昌矿业武庄铁矿正义之窗9求助！求助！我们农民工辛苦挣了一年钱！到了年头最基本的工资都拿不到！要工资要了五个月了！找政府！政府说管不了！找龙成集团许昌铁矿！他们说没有钱！我农民工工资就这样没有了着落了！可怜我农民工！希望有能力人事和媒体给帮帮忙为我们作主！求转发！扩散！大家帮帮我们可怜的农民工          我们农民工在河南许昌县苏桥镇！武庄铁矿干了半年活！临近年关了！二百多工人的工资一分钱没有！矿方不给工头结账！工人问工头要工资！工头吓跑了！而矿方现在不管工人了！ 工人现在没有吃的！没有喝的！还拿不到基本的血汗钱！希望朋友和媒体给我们农民工伸张正义！＊［工人］2015.1.22 湖北 宜昌市 猇亭区 华润电厂*********狼了这是个什么世道！宜昌猇亭华润电厂大门口农民工拿起横幅讨血汗钱 还有人扬言要拿钱请人殴打这些农民工 警察来了不帮农民工反而强行收走横幅 请社会各界人士关注 农民工幸苦一年很不容易。竟然还有这样黑心的老板 让人心寒！农民工不容易 拿个工资怎么就这么难 都说社会是公平的 但它体现在哪里呢。警察都帮着老板 这公道在哪？＊［工人］2015.1.22 四川 成都市 双流县 益端鞋业有限公司何奇晋希望有关部门解决这事 农民工工资不能拖欠哦 年底了 工人们都等着钱回家与家人团聚。＊［工人］2015.1.22 四川省 绵阳市 游仙区 游仙镇 石垭村统建房BingBange又是年终农民工讨薪！横幅都拉到政府门口了 该给个说法吧！＊［工人］2015.1.22 河南 平顶山市 鲁山县 圣光医用制品有限公司平常心828408（横幅：变相裁员拒不赔偿）内地老板仗着与政府管员有关系 漠视弱势群体的利益 曾几何时 在沿海一带也是经常上演 只是到年关了 叫人怎么活呀！蝶雨829 （圣光）圣光还我血汗钱1、平顶山神行保健科技有限公司迄今为止 公司已拖欠2个月工资没有发放（2014年11月和2014年12月份工资两个月 公司规定 工资应于15日前发放上一月的工资）。2、平顶山神行保健科技有限公司存在变相裁人 但平顶山神行保健科技有限公司未按照国家相关的法律法规给予陪偿 2015年1月17日（周六）由各部门领导口头通知（没有正式的文件）大部分办公室职员即日起正式放假3个月 经1月20日我们到鲁山劳动局提出请求劳动仲裁后 公司才临时通知放假期间公司给出的薪资待遇为：农村户口110元/月、非农村户口300/月的补助。此举已严重违反国家相关法律。1月20日中午从劳动局回公司后 我等部分员工才收到领导转发的短信及口头通知 短信内容为：“转达人事部关于人员淡季放假安排及辞工结算事项 现因业务淡期 统一长假从1月16日至4月16 期间公司按照劳动部门规定发放最低生活费 若因个人原因在1月20日至21日两日内提交辞工申请的 1月份工资按全月工资发放 23号起行政部统一收缴桌椅、电脑等公司资源 以上具体安排以人事部文件为准。”3. 公司已数月未曾为员工缴纳统筹 相关保险等 已严重违反相关法律法规。＊［工人］2015.1.22 福建 漳州市DP32Hazel瑄回家路上眼都看呆了现场群情激愤都快打起来了[发抖]110们都把道路封锁起来了车辆无法进入.福海阳光现场示威口号震耳欲聋。＊［工人］2015.1.22 湖北省 宜昌市 夷陵区 鸦鹊岭镇 罗汉生态红提休闲庄园暮雨18宜昌鸦鹊岭政府 农民工讨薪！＊［工人］2015.1.22 福建省 漳州市 漳浦县 杜浔镇学超Ren（陈乔华曾爱清还我血汗钱）农民工堵路讨债。杜浔 ＊［工人］2015.1.22 陕西 西安市 未央区政府不转身已陌路中央不是说了嘛！必须保证农民工工资不拖欠 可是这是为什么呢？？？＊［工人］2015.1.22 海南 三亚市 龙泉谷·三亚的山（中度）golf小青青快过年了！大家辛辛苦苦忙活了一年容易吗 还拖欠农民工的血汗钱golf韩小颜快过年了 坑爹的房地商们拖欠农民工的务工费 拦路要款 希望他们顺利拿到自己的辛苦费开心回家过年＊［工人］2015.1.22 河南省 新乡市 获嘉县 太山镇 辛章村说说新乡事儿亲们 金穗大道公园南门农民堵路中 请绕行瑾柘人民公园南门堵路了 请绕行！＊［工人］2015.1.22 湖北 咸宁市 崇阳县 兴民钢圈hubeixiaohuang咸宁市崇阳县兴民钢圈欠建厂房的农民工30多人的工资不给 有政府袒护 县政府领导拿烟灰缸砸农民工 警察也拿警棍打农民打农民 ＊［工人］2015.1.22 河北省 邢台市 清河县牛逼的King拖欠农民工工资。Gareence农民工的工资不可拖欠 都交通堵塞惹！＊［工人］2015.1.22 江苏省 徐州市 铜山区 马坡镇jh**********这就是江苏省徐州市铜山区马坡镇的中国人民警察不为人民的哦！农民工要血汗钱 他们在前面拦住不让要。警察现在就是以前国党的二狗子狗汗奸。还说我们要钱是围法的 我们不这个工地上四个月没拿一分钱。政府公安都是要喝我们建筑工人的血哦！请有关部门帮帮我们哦！不会让我们真的要去跳楼吧＊［工人］2015.1.22 广东 广州市 佳兆业城市广场刚被T了佳兆业 城市广场项目 工人讨薪堵路＊［工人］2015.1.22 江西 南昌市倔强的思彤小姐往丰城去的那条路上 堵死 又是老板拖欠农民工工钱 导致做出这么过激的事情 政府部门年年讲着要为百姓解决这类的事情 可有时候就是山高皇帝远啊＊［工人］2015.1.22 广东 深圳市 深中润集团庚戌年偶遇的抗议事件 希望他们可以过个好年 ＊［工人］2015.1.22 贵州省 遵义市 遵义县 南白镇小汤圆love源子农民工讨薪＊［工人］2015.1.22 陕西 榆林市 子洲县 永兴煤矿用户**********子洲县永兴煤矿拖欠农民工资一年多 多次索要受到老板雇佣黑社会组织来矿威胁 无奈多次去县政府给予帮助 却操蛋的奇葩 我们解决不了来到榆林市政府门口 又一次遭到门卫镇压 说是影响市容 最后说让我们去信访局 可来到信访局 六点了没人来解决此事 这难道是我们老百姓心中的政府 痛哉 哀哉？＊［工人］2015.1.22 安徽省 安庆市 望江县政府清道夫2012-2#安徽望江县群众路线搞得好#驰名中外的办公楼＿赛白宫（望江县委县政府）门口经常聚集大批警察 他们对付的就是讨要工资的农民工。＊［工人］2015.1.22 黑龙江 齐齐哈尔市 富拉尔基区 天河湾讨薪难难北京上访。齐齐哈尔富拉尔基天河湾小区 农民工艰难讨薪 处处受限制 O微博视频李晶ld去北京告状 老百姓容易吗 农民工的血汗钱都不给。黑龙江的农民工去北京找开发商要钱。＊［工人］2015.1.22 云南 昆明市 海伦国际__虢景荣昆明广福路被堵 海伦国际工人游街闹事 和警察打起来了。起大风了吗海伦国际。农民工讨薪却没有政府部门的人来管.后来。来了一帮警察和几个协警。一来就打这些.讨要工资的农民工。这些政府太污了。大家帮忙转起来吧！谢谢瓜尔佳茉雅奇这些农民工太可怜啦 海伦国际不付工钱85H小警广福路发生堵路事件。 O微博视频找片和谐广福路上、全是海伦国际的讨薪农民工！漠视********伤不起的讨薪族 伤不起的广福路 伤不起年代 除了看看热闹外也无能为力＊［工人］2015.1.22 海南 儋州市 东风派出所勤奋的紫衣大侠海南省儋州市农民工讨薪 谁知儋州市政府和欠薪老板钟丽新同流合污 派警察镇压殴打农民工 并抢夺农民工手里的资料 企图毁灭证据 逃避欠款。其中儋州市东风派出所所谓的副所长 警员编号PC140479 更是牛逼哄哄 为钟丽新出头。可怜的农民工一天讨薪未果 儋州市政府不理不睬 只能睡在马路边。＊［工人］2015.1.22 陕西 安康市 宁陕县 宁陕新天地／邦柯建筑劳务有限公司任国栋爱娇娇宁陕新天地邦柯劳务公司拖欠民工工资。找政府处理然而一拖在拖整整拖了半年。现在过年工人都在宁陕县政府肯求解决。但是县政府却一推在推 现在民工也饭都吃不起住不起。老人喊天理何在。 ＊［工人］2015.1.22 北京市 通州区 辉煌时代家具有限公司张咪-足迹北京市通州区马驹桥小周易村 辉煌时代家具有限公司 拖欠工人四个月工资不发。求广朋友用你们万能的微博朋友圈往死里刷。谢谢。拜托＊［工人］2015.1.22 湖北 荆州市 荆州区 弥市大桥Diligent_梅子弥市大桥今天又被堵了 昨天也进行了这样的事情！农民工拿不到工钱回家过年 无人管他们！为了生计 他们不得不采取这样的做法！可是也因为这样 交通瘫痪 这样又害了多少有急事的人们！快过年了 希望这件事情能够尽快解决 农民工们能回家过年＊［工人］2015.1.22 河北 邯郸市 武安市 运丰冶金工业有限公司512佳珊河北省武安市矿山镇崔石门村村南 《运丰钢铁冶金有限公司》。 老板崔运生 拖欠全公司1千名员工8个多月工资不发 还不让员工辞职。 电话投诉石家庄 石家庄推给邯郸 邯郸推给武安 武安推给矿山镇。 员工一年辛辛苦苦的血汗钱到头来不给 难道非得捅到中央你们才管吗? 望广大群众看到此贴的转起来 武安苦命人河北省武安市运丰员工上访讨要七个月工资！＊［工人］2015.1.22 河北 唐山市 开滦（集团）有限责任公司唐老呔儿实时报道 开滦工人又开始集结 讨要辛苦劳作应得的工资！条幅打出来了 还我血汗钱！＊［工人］2015.1.22 （江苏省 无锡市 江阴市 祝塘镇）用户r6hejzji39祝塘某服装厂拖欠员工工资 老板不发工资 还好意思报警。又罢工了 老板又不发 老是拖欠员工工资 真是不想给他干活了 真不要脸。＊［工人］2015.1.22 安徽 合肥市 安徽广电草根合肥年关了 安徽广电居然也被农民工拉横幅讨薪了VIA@雨甜-oo＊［工人］2015.1.22 云南 文山市 金昆房地产八次以后 （农）农民工要工钱来交通宾馆堵路了。据了解是农民工来早工钱。是云龙商场工地那里的工人。文山村民 金昆公司风光不再 危机四伏！＊［医护］2015.1.22 江苏省 南通市 如东县意料之外的浪漫情书（横幅：回归公立医院；恢复事业单位编制）江苏省如东县乡镇卫生人员请愿县政府＊［农民］2015.1.22 广东省 汕头市 潮阳区 西胪镇 西一村MIM2A传说中的汕头市潮阳区西胪镇人民与开发商 与村官示威的一小场景。远超过80亩的农田变建设用地 既然合法 那么阻止上访 及电台报道又是闹什么？可怜的人民。＊［农民］2015.1.22 山西省 太原市 万柏林区 长风街道 小王村西瓜是草莓味2小王村村民注意。大家要团结。反腐败坚持抵制腐败现象。原本的公园现在居然要盖小区。大家好好想想。小王村腐败现象已经这么严重。大家团结起来。求转发你好逗z小王村村民你们都是好样的 不能在让那些贪官们逍遥法外了。-苗德强求转发：山西省太原市南内环小王村官员贪污。腐败严重。小王村村民要团结。反腐败斗争要坚持。官员官官相互 中饱私囊 层层勾结 祸害村民利益。破坏村民安居乐业生活。＊［农民］2015.1.22 河南 郑州市 经开区 九龙镇 席庄村_方枪枪没有小红花四港联动大道九龙镇的十字路口又发生村民堵路事件 以前因为村民过马路出交通事故多次堵路 这次好像是因为路口红绿灯不亮 村民想修红绿灯又来堵路…走这条路的司机也经常闯红绿灯 村民安全出行也是一大问题。真不知道到底是谁的责任文艺范chuan目前四港联动大道几辆货车横在路中间 堵路了 过不去 我在四港联动大道郑尚线嘻嘻呵呵2 （我反映）我反映的是有关交通安全的问题 车祸猛于虎 人命重如天。在四港联动大道与经开区九龙镇席庄村处的十字路口 经常发生车祸 这个路口是附近村民赶集的必要通道 人流量很大 可是这个路口的交通信号灯形同虚设 南北过往的车辆根本就不遵守交通规则 多数车辆闯红灯 而且速度也很快 给当地的村民生产生活带来了极大的安全隐患 恳请 领导关注一下 解决我们出行的后顾之忧。＊［农民］2015.1.22 四川省 内江市 东兴区人生若只如初见cheng大清早出门就遇到这种事 一大群人横拦在马路中间 不让任何车辆过 看到他们横幅上说“贪官强卖林”什么的 大帮人来拦路一女的还和过路一司机打起了 车上人都议论 要讨公道去区政府 市政府嘛 拦路拦我们咋子都不晓得 真的是！堵了我半小时！内江东兴区 修高铁站这边＊［农民］2015.1.22 山西 长治县 小河南村婷子tiing小河南村的老百姓维护自身合法权益从乡到县再到市投告无门 政府一再推脱不予以一个说法 被逼无奈之下跪求在市政府大门前 一个个村民看着眼前树立的大石碑上的“为人民服务”心里是何感想？可悲可怜可怒可恨 这就是所谓的伟大的中华民族耻辱＊［农民］2015.1.22 安徽 合肥市李小喂LIVE你们tmd除了腐败镇压你们还会什么？无知狗 。开发商和农民发生土地纠纷 开发商不解决。政府出特警镇压解决。腐败的政府 痛心＊［拆迁户］2015.1.22 湖北 武汉市 汉阳区 知音桥疯叶-秋诗一个爹爹因为政府强拆被打伤 一群爹爹婆婆上知音桥开始堵桥！说好的和谐文明城市呢？特警和防爆队都出动了！海堂花不会自己开一些老人把路堵了抗议 武汉市江汉二桥桥头阿狸狸狸de桃子知音桥好可怕。第一次碰到这样的情况 一群爹爹婆婆睡在路中间 其中一位婆婆还给我们看床上那个受伤人的断腿 整个王家湾都被堵了 车进不去 出不来 之后走回来的时候看到好多特警 不知道后来处理的怎样Bordeaux吴知音桥废了 搞不清白带闹么事 一群爹爹婆婆带中间堵马路……就算有么事不平的也不能这样搞撒 害人 特警都来了。。。small_魔_girl_大家不要走知音桥～维权的婆婆们把床抬到桥上来了对不起这名字 （二桥）二桥又有人静坐堵路了。不要命了 吊着水也躺床上上来了。＊［商户］2015.1.22 湖北 武汉市 江岸区 幸福时代幸福里商业街乐熙妈妈武汉市江岸区百步亭幸福时代商业街黑心开发商跟警察流氓勾结对付业主商户 停水停电 天理何在…帮忙关注＊［业主］2015.1.22 黑龙江 哈尔滨市 地一大道香港城（人和四期）-__天道酬勤__-在习主席领导的年代 解决问题得下跪。黑龙江哈尔滨 260多名黑龙江的老百姓给您再次下跪 请求市委领导出面解决人和四期香港城欺骗1300多户业主上亿人民币一事。还老百姓一辈子的血汗钱 恳请市委有领导站出来 为老百姓主持公道！＊［业主］2015.1.22 辽宁 朝阳市 圣煜房产陈丽斌斌辽宁省朝阳市环保局和圣煜房产公司在没有预售许可证情况下组织团购卖房438户 开发商预先使用团购预付款1亿以上近三年之久 现既没按合同13年底交工 也没按合同承诺团购户多层房而是高层 多次找政府协商 结果只高层 开发商没钱！可怜的百姓们只能踏上访之路了！＊［业主］2015.1.22 贵州 贵阳市野猫瞳房子什么时候才能见到你 无良房开经济房修成烂尾楼 业主要求政府给说法。＊［业主］2015.1.22 黑龙江 哈尔滨市 星光耀广场蝙蝠侠的小超人曾经万众瞩目的星光耀 如今面临如此局面你们是何感想@哈尔滨星光耀广场官方微博？你们欺骗业主购房时 是怎么忍心说出那些谎话的？业主维权时 又是怎么忍心找社会人威胁恐吓的？你们没有父母？没有儿女？动手打人 难道没人管了吗？习大大当道 你们如此放肆 勾结官员 收买媒体！不会有好下场的！＊［死者家属］2015.1.22 广东 茂名市中医院茂名娱乐网[今日关注]网友爆料称 他今天上午去了趟中医院 发现门口100来个防爆警察 后来听中医院里面的人说刚才有大批人围堵医院 说是医院治死人了 家属还在门口烧香。现在的医院是怎么了？＊［退伍军人］2015.1.22 广东 阳江市政府看二看 （市政）市政府又无知发生咪事 好多人。边个来讲解吓。我爱龙津路女生 不是讨薪 是对越作战复退军人要求提高保障待遇＊［退伍军人］2015.1.22 山东 聊城市政府wg峰哥888 （主题：）主题：市政府门口热闹了 莘县和临清的自卫站老兵在市政府门口上访 要求享受同等待遇 支持＊［退伍军人、军属］2015.1.22 河北省 张家口市 赤城县厾亓籁籁河北省张家口市赤诚县人民政府欺骗退休军人即家属 退伍军人即家属要求政府兑现承诺 家属长跪政府门口 政府官员无动于衷 县委书记更是坐在车上始终不下车！求好友们转发！用户**********河北张家口市赤城县 2013年复原军人因安置问题不明 面见政府 答案含糊不清 推推拖拖。政府门前军属长跪不起 书记置之不理 这就是人民政府 这就是党领导下的班子 这就是保家卫国 复原军人应有的待遇 寒心啊。小小＊［投资人］2015.1.22 四川省 遂宁市 射洪县 铭亿融资理财信息咨询有限公司供水小唐勿有贪念 射洪县投资公司跑路了 老百姓讨说法堵路了 唉 太坏了慧质岚馨1025特警出动了……搞凶了……勤奋的罗luo （堵路）堵路了国色酒香 （铭亿）铭亿又遭了 罢路 强大的可有？＊［投资人］2015.1.22 湖南 长沙市 博沣资产管理有限公司Q天山飞雪遭遇工商银行理财产品骗局的受害人 今天聚集到湖南省委上访维权 希望事件能得到妥善解决！＊［投资人］2015.1.22 河南 开封市 北京大汗天下传媒有限公司开封分公司K-K-O又见开封堵路 原来是大汉天下也倒了~哈哈哈 你投资拍个《洋妞到我家》也没见你多牛逼~哎~切莫盲目贪图高息啊~非池中81 （汉兴）汉兴路又堵路了 大家绕行吧 又堵路了 人山人海啊 啥都过不去房倒屋塌中 :大汗天下门口 好像又是投资公司。据说这都是大客户 起步十万。＊2015.1.22 河南 郑州市 紫辰路／紫东路oO鄭州龍Oo紫辰路紫东路口闹事堵路了 不清楚原因林小飞_紫辰路与紫东路被些刁民堵了交通严重瘫痪 ＊2015.1.22 江西省 景德镇市 浮梁县 寿安镇 仙槎村 窑坞煤矿绾君歆1618仙槎煤矿门口拦路。公交车都堵了2辆 后面跟的打的个走涌山绕的一圈走噢＊2015.1.22 湖北省 黄冈市 麻城市 中一镇政府QQ*******群众在中一镇政府门口上纺＊2015.1.22 河南 新乡市兔宝宝的夏小天市级执法人员常宝柱与新乡宾馆陈红串通一气 污蔑百姓 扭曲事实 颠倒黑白 强行将老百姓连拖带拽拉进其执法车内进行殴打 有违国法 天理难容 后以办完事为由请客吃饭 目无王法 天理难容。还我公道！跪求扩散！！！我们希望你动一下手指。帮我们转发一下。＊2015.1.22 （湖南 长沙市）羊晓小羊在马路中间排排站还拉起了横幅 这是怎么了？＊2015.1.22 上海市 徐汇区政府百合奇琪徐汇区区政府门口是怎么了？会有新闻吗?＊2015.1.22 上海阳晨排水运营有限公司闪闪发光的女神金（横幅：欺诈合同 违规违法停水停电）一大早上班路上看见的 在抗议龙华排水厂 群众在排排坐吃包子。啥情况这是？？龙漕路附近吧＊2015.1.22 河南 商丘市 永城市委用第六套广播体操轻松击败你永城市委门口。好多人不知道干嘛的。＊2015.1.22 湖南 衡阳市政府胡-歌V又见上访＊2015.1.22 贵州 遵义市 仁怀市谭老大想去伊瓜苏出门遇到喊冤封路 特警镇压 太暴力 冒死偷拍我想我能从事记者行业！"|http://newsworthknowingcn.blogspot.com/2015/01/2015-01-22.html|2015-01-24
其他媒体|1750769238|163|网易文化论坛-活动专区|ZHO|2015-04-13 23:17:01|我的首台双系统平板 - 蓝魔i11pro体验|两周前我收到了蓝魔i11pro平板电脑 在这半个月的时间里 我充分地体验并观察这款为数不多的双系统平板 并没有急于分享也是我一贯的态度。回想去年9月份的发布会至今 蓝魔与因特尔 比亚迪合作推出了包括i7s i9s i10s在内的一系列产品。一转眼i11pro也到来 它给我印象最深的两点就是：①双系统的实用 ②超大尺寸的震撼。使用中也总结出存在的问题 就听我简单快速地分享之。        ★包装简约中肯                     传统开箱就不做重点 一笔带过也就是了。我总共收到两个独立包装 分别是机器和订制键盘。配置采用阿童木凌动处理器（atom z3735F） 10.6寸1080P 2G内存 32G eMMc 还有售后信息都写在背面。因为10.6尺寸并不常见 键盘并不能与市面10.1平板通用。        ★外观漂亮 配件不够丰富                  其他附件并不多 包含数据线 充电器 说明书 合格证。并没有otg线 这对日后使用造成不小的麻烦（后面详细说）。                  正面1080P IPS屏非常震撼 相比1920 x 1200 的10.1寸平板更宽一些 有着不错的观影效果。简洁为主 并没有什么花哨的装饰。                  平板右侧有一个圆形虚拟键 这实际上是WIN8.1系统下的HOME键。我以前用的WIN平板多是微软徽标 并且出现在下边框 所以刚开始有些奇怪。在Andriod系统中这个虚拟键没有实际作用。                另一个问题也是比较突出的 唯一一个Micro usb既要负责数据传输 也要负责充电 不是很方便。标准usb接口的缺失 意味着同时使用优盘 蓝牙设备（鼠标 手柄等）产生矛盾 只好添加HUB来缓解一下。                  相比前作之一的i9s i11pro在工艺上有所变化 正面依然采用钢化玻璃 后壳则改为一体成型铝合金材质 并且加入喷砂工艺。这些改变很难说孰优孰劣 喜好也因人而异。                  机身左侧排列两个实体键 启动键和音量键 并无什么特别之处。反馈明确 键程舒适。一圈金属包边 严丝合缝。2.5D圆角提升外观的立体感。                     前文提及到 10.6寸并不多见 键盘也需要特殊订制。Docking触点并无特别 但是其两侧的固定卡扣略有不同。现在还不能确定标配是否一定送键盘 若不送可不能随意选择10.1寸的磁吸键盘对付哦。        ★功能强大的双系统                  蓝魔最近的系列产品中 以pro后缀的都是双系统。这里面包含已经被玩烂的安卓系统（Andriod4.4版本） 和刚兴起不太久的微软系统（Windows8.1）。前者侧重娱乐 后者注重商务。目前为止i11pro还不支持热切换 开机时才能选择何种系统。启动速度很快 这点不错。                  别怪我偏心 一年前我就不太专注安卓平板了 这和手机尺寸日益扩大化 手机系统更新换代速度 优秀地订制程度有关。所以我就先从Win8.1说起。相信Metro桌面大家都非常熟悉啦 贴近上下左右四个边框向中间滑动的手势 对于初学者还是相当有吸引力的。注册并登陆微软系统 实现更多复杂的功能 如：note 微软市场 必应系列app等。或者直接采用本地离线账户 但不推荐。App的种类繁多 但不符合国人的口味 感觉有点杂乱。                  而切换传统桌面后就和笔记本无异了。你会发现程序运行方式 操作手法都很熟悉。在这种状态下推荐使用蓝牙鼠标 更加舒适。键盘输入在办公室得心应手。软件兼容性很强 不会出现当初xp跃进Vista时出现多程序不能运行的现象。我的i11pro为32GB版本 均等的双分区 分别安放两个系统。但在各自的系统时不能写入另一个分区（虽安装特定软件后仅可以交叉读取 但也不是很方便）。容量就不太够用 WIN8.1中尤为明显。最好的办法是通过底侧的TF卡槽扩展作为仓库盘。考虑到32G和64G只差100元 推荐后者才是王道。              出厂系统已激活 但是没有赠送office激活码 所以我需要通过一些软件破解一下 一般在网上下的win8.1系统内都有 我就是从装win8.1的台式机上拷贝下来哒。有时候外出需要晚上赶稿件 带笔记本又不方便就用它。                     无聊时也可以打点游戏 一般的大型3D游戏都能成功运行 测试了使命召唤5-世界之战 720P下比较勉强 激励场景略有卡顿 目测帧数20左右。尘埃2不是fps类型 视角转换较小 所以流畅度明显高于前者。整体体验下来有较高体验水平。通过大型游戏也能大致评估i11pro的性能 对付其他一般的办公软件 甚至叫专业作图软件都能轻松应对。                     再来体验安卓4.4操作系统 这个系统相对简单 也被大家熟知。键盘除了体现输入优势外 几乎也就当个支架 所以更多时候是拿下来捧着玩。X86构架 64bit的z3735F相比传统ARM（如：rk3288 A80）性能提升太明显 第七代Intel Graphics芯拥有强大的图像处理 使用时感觉极为流畅。                  默认谷歌浏览器 字体 字号我认为比WIN系统的漂亮清楚。同样支持多页面选项卡切换 但不能像win8.1里ie11那样同时运行。                     大屏下最舒适的就是观看图片和电影 这是我第一次使用10.6寸的平板电脑 比14.1寸小不了多少 但是轻便许多。质量稍重 不适合长久握持。1080P显示分辨不算视网膜 细腻程度也不错。IPS屏178°广视角 令人满意。期待加大内存 提高称4k屏幕。                  开启intel独有的视频优化 解码更加轻松流畅。                  双系统有个非常实用的用法 就是如果WIN系统搞崩溃了 可以在Andriod里恢复WIN系统 对于不会重装系统的小白太方便了。                  自带的谷歌软件市场一般 登录谷歌账户之后可以下载些app。但是我还是习惯用豌豆荚和当乐游戏中心。里面超多免费 破解游戏。因为配置过于强大 安卓平台的游戏还没有不能玩的。        【总结】        这么多天使用下来基本满意 百分制衡量的话我会给85分。外观 性能 尺寸 双系统是我较为满意的。WIN系统下字体很小 虽然可以通过修改字号 调低分辨率等方法有所改变 但是终究在办公的时候稍显吃力。最后如果能在后期加上标准usb 更改为DC充电器的方式 加大内存 提高到4k分辨率 将会是一款完美之作。|http://club.tech.163.com/bbs/mobile_activ/528797808.html|2015-04-13
其他媒体|1773056041|sohu|大话it|ZHO|2015-04-27 21:14:02|直击上海车展 比亚迪新能源车阵容新员解析|新泽西州   性别:未公开 所在地:未知 社区生日:未知   发帖总数:0  精华帖数:0 声望魅力:0 积分:0     送礼物 留言 关注 加好友   楼主   昨天刚看完车展 今年比亚迪展台展出的全部都是新能源车 难怪自称为新能源车的领导者 还没见哪个车企在新能源车这块儿做的这么投入 做的这么专业。一直对比亚迪的新能源车比较关注 尤其是比亚迪秦 油耗低、外观漂亮回头率高 空间大 混合动力强劲 完全颠覆了我对传统汽车的认识 从那时候起我就默默的变成了一名小迪粉儿。这次逛车展看到比亚迪又发布了两辆新能源车 一个是“宋” 一个是”元“ 这是两款混合动力的SUV 这回比亚迪的新能源车的阵容又壮大了。“宋“是一款三擎四驱双模SUV 百公里加速时间在5秒以内 这动力性系统确实够牛的。  宋的外观与以往比亚迪车型的外观不太一样 运用全新的设计语言 前脸采用X型的装饰板 配以犀利的前大灯 整个车头看上去非常有冲击力 运动感十足。车身前后logo下都配有前摄像头 这个倒是挺实用的。车身的颜色上下不一样 车顶有行李架 车身侧面腰线上扬 使整体外观看上去都动感十足。不过比亚迪的车身尺寸比唐略小一些 4565*1830*1720mm的车身尺寸 2660mm的轴距 还是符合它是一款中型SUV的定位的。轮毂造型别致 米其林LATITUDE轮胎挺厚道。内饰方面 全黑的内饰配以仿实木花纹的装饰板 整体感觉比较上档次 仪表盘虽说不是全液晶的 不过该显示的读数还是都有的 也比较直观。方向盘的握感也比较好 液晶显示屏、PM2.5绿净都有 座椅的舒适性不错 空间比我想象中的要大。大天窗 各功能键的布局合理 总得来说宋的内饰设计还是相当人性化的。            接下来再聊聊元 “元“是一款小型SUV 长宽高分别为4320/1765/1650mm 轴距2520mm 尺寸上比宋略小 不过外观同样是走运动路线。不管是黑白蓝的配色 还是线条感十足的外观设计 再加上犀利的大灯 元给我的事一种小硬汉的感觉 多幅式轮毂更是点睛之笔。 车尾的设计给我留下印象挺深刻的 外挂式备胎采用类似于旋转风车的设计 门把手隐藏在车尾大灯的位置 这样的设计刚开始觉得挺不可思议 不过看过车你就知道 绝对没有突兀之感。“元”的动力系统由一台1.5L的自然吸气发动机 还有两台电动机组成 同样的四轮驱动。纯油的情况下 1.5L的动力对于元的车重来说完全算得上动力充沛。在纯电动模式下 最大续航里程同样可以达到70公里。看车的时候没拍到内饰 因为不让进去 不过就在外面看 元的内饰材质和做工还是挺细致的 该有的功能也都有。        这次车展比亚迪携旗下的唐、宋、元、商 纯电动出租车e5、纯电动物流车T3等等新能源车参展 比亚迪的新能源车的队伍确实挺强大。比亚迪还发布了新能源车“7+4”全市场战略布局 看来未来比亚迪的新能源车的阵容还会不断壮大。              只看楼主    回复     举报  发表于 15-04-27  20:06:30   新泽西州的签名档|http://club.it.sohu.com/it/thread/35k3ulmxhg9|2015-04-27
其他媒体|1805361194|hexun|滚动新闻 > 全部新闻|ZHO|2015-05-17 20:11:02|优惠靠诚心：2014起亚k3多少钱 2014起亚k3试驾|　　店内促销火爆进行 起亚k3最高优惠3万元 并有全车精品2.5万装饰赠送 目前店内有现车充足 颜色齐全 对该车感兴趣的朋友可致电经销商详询 销售热线：010-59******-*******3930李经理　　起亚K3最新报价表车型(北京报价)指导价(万)4s店价格(万)价格变化(万)备注1.6L 手动GL2014款10.287.283现车1.6L 自动GL2014款11.288.283现车1.6L 手动GLS2014款11.488.483现车1.6L 自动GLS2014款12.489.483现车1.6L 自动DLX2014款13.1810.183现车1.6L 自动Premium2014款14.3811.383现车1.8L 自动Premium2014款14.9811.983现车销售热线：010-59******-*******3930李经理　　『起亚K320141.6L 手动GL』　　外观上 2014款K3秉承“Design KIA”设计理念精髓 在车身前脸和尾部均有全新呈现。前脸全新的前中网颜色 使得虎啸式家族脸谱视觉感受更为动感大气且引人注目。　　内饰方面 K3在中控面板等部位进行了软性涂装 并且在空调按钮处增加了镀铬装饰和旋钮形状的改善 质感升级带来细腻的触感 让驾驶者身心愉悦。K3动力系统搭载1.6L和1.8L发动机 并且配备6速手动或者6速手自一体变速箱。　　编辑点评：起亚K3外观时尚动感 内饰中控台按钮简洁 功能配置齐全 车内空间表现不错。起亚K3是与北京现代朗动同平台的一款紧凑型轿车 该车外观时尚美观 拥有优美的线条 内饰具有科技感 很强的运动风格 同时该车采用了1.6L和1.8L两种排量发动机可供选择。　　五星级诚信企业　　更多详情可致电经销商：010-59******-*******3930李经理　　是否现车：现车齐全　　经销商名称：北京隆翔汽车销售服务有限公司　　经销商地址：北京市朝阳区北五环外立水桥69号。　　《北京地铁五号线天通苑站下车往北200米》　　下车电话联系有专车接送。　　以上信息仅供参考 具体优惠信息以到店核算为主。　　如系本站原创文章 转载请注明出处：汽车中国。（责任编辑：HN666）|http://auto.hexun.com/2015-05-17/175884353.html|2015-05-17
其他媒体|1864308618|zhidao_baidu|生活|ZHO|2015-06-20 21:44:01|东风悦达起亚k3是仿美车型|来自：手机知道生活|http://zhidao.baidu.com/question/177520375570868724.html?entry=qb_browse_default|2015-06-20
其他媒体|1897548534|hefei|合肥专区|ZHO|2015-07-10 00:03:02|2015年甘肃省一万名考试题 答案《★７********★》|"2015年甘肃省一万名考试题 答案《★７********★》  2015年甘肃省一万名考试 答案【通过率100%卡卡客服Ｑ７********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年甘肃省一万名考试真题答案-2015年甘肃省一万名试题及 答案-2015年甘肃省一万名考试时间-2015年甘肃省一万名进村进社考试科目-2015年甘肃省一万名考试大纲-2015年甘肃省一万名考前答案-2015年甘肃省一万名答案【Q７********包过】-2015年甘肃省一万名考试资料【Q７********包过】-2015年甘肃省一万名复习资料-2015年甘肃省一万名考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级甘肃省一万名著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年甘肃省一万名考试 答案=７********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级甘肃省一万名考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年甘肃省一万名考试 答案 试题 真题 时间 科目〃Ｑ７******** ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年甘肃省一万名考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年甘肃省一万名考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案７********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=７********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级甘肃省一万名考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=７********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级甘肃省一万名考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级甘肃省一万名考试 答案=７********.祈福2015年甘肃省一万名进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年甘肃省一万名考试 考式 答案=７********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年甘肃省一万名考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=７********人时简累 会受苦 正高级高级甘肃省一万名考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=７********.祈福2015年甘肃省一万名考试 考式 答案=７********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级甘肃省一万名考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=７********.祈福2015年甘肃省一万名考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=７******** ^1 q) ~# t: {/ h/ J【=７********.祈福2015年甘肃省一万名考试 考式 答案=７******** W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年甘肃省一万名考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. ７********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年甘肃省一万名考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=７********.祈福2015年甘肃省一万名考试 考式 答案=７********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级甘肃省一万名考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=７********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级甘肃省一万名答案【Q７********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级甘肃省一万名考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=７******** 2015年甘肃省一万名考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年甘肃省一万名考试 考式 答案=７********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年甘肃省一万名考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=７******** 2015年甘肃省一万名考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级甘肃省一万名考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W７********=７******** 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^７********_100%】哪个2015年甘肃省一万名考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=７********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年甘肃省一万名考试 考式 答案=７********.+ F; ~ C( X7 G$ ?$ I祈福2015年甘肃省一万名考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年甘肃省一万名考试 考式 答案=７********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级甘肃省一万名答案【Q７********】9 I' [+ v* p3 m' Q=７********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级甘肃省一万名 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年甘肃省一万名考试 考式 答案=７********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级甘肃省一万名考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=７********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年甘肃省一万名考试 考式 答案=７********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级甘肃省一万名考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=７********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”７********.祈福2015年甘肃省一万名考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级甘肃省一万名考试/ J7 J' y9 ]5 c5 w; D答案=７********.祈福2015年甘肃省一万名考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级甘肃省一万名考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年甘肃省一万名考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案７********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=７********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年甘肃省一万名考试 答案Ｑ７********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15326119&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-07-10
其他媒体|1897604657|hefei|合肥专区|ZHO|2015-07-10 00:42:01|2015年甘肃省一万名考试题 答案《★280119７75★》考后付|"2015年甘肃省一万名考试题 答案《★280119７75★》考后付  2015年甘肃省一万名考试 答案【通过率100%卡卡客服Ｑ280119７75包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年甘肃省一万名考试真题答案-2015年甘肃省一万名试题及 答案-2015年甘肃省一万名考试时间-2015年甘肃省一万名进村进社考试科目-2015年甘肃省一万名考试大纲-2015年甘肃省一万名考前答案-2015年甘肃省一万名答案【Q280119７75包过】-2015年甘肃省一万名考试资料【Q280119７75包过】-2015年甘肃省一万名复习资料-2015年甘肃省一万名考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级甘肃省一万名著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年甘肃省一万名考试 答案=280119７75- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级甘肃省一万名考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年甘肃省一万名考试 答案 试题 真题 时间 科目〃Ｑ280119７75 ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年甘肃省一万名考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年甘肃省一万名考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案280119７75.祈福2015年内蒙古会计从业资ac格考试 考式 答案=280119７75+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级甘肃省一万名考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=280119７75人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级甘肃省一万名考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级甘肃省一万名考试 答案=280119７75.祈福2015年甘肃省一万名进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年甘肃省一万名考试 考式 答案=280119７75.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年甘肃省一万名考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=280119７75人时简累 会受苦 正高级高级甘肃省一万名考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=280119７75.祈福2015年甘肃省一万名考试 考式 答案=280119７75人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级甘肃省一万名考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=280119７75.祈福2015年甘肃省一万名考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=280119７75 ^1 q) ~# t: {/ h/ J【=280119７75.祈福2015年甘肃省一万名考试 考式 答案=280119７75 W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年甘肃省一万名考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. 280119７75[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年甘肃省一万名考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=280119７75.祈福2015年甘肃省一万名考试 考式 答案=280119７75人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级甘肃省一万名考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=280119７75_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级甘肃省一万名答案【Q280119７75】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级甘肃省一万名考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=280119７75 2015年甘肃省一万名考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年甘肃省一万名考试 考式 答案=280119７75.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年甘肃省一万名考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=280119７75 2015年甘肃省一万名考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级甘肃省一万名考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W280119７75=280119７75 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^280119７75_100%】哪个2015年甘肃省一万名考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=280119７75人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年甘肃省一万名考试 考式 答案=280119７75.+ F; ~ C( X7 G$ ?$ I祈福2015年甘肃省一万名考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年甘肃省一万名考试 考式 答案=280119７75.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级甘肃省一万名答案【Q280119７75】9 I' [+ v* p3 m' Q=280119７75⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级甘肃省一万名 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年甘肃省一万名考试 考式 答案=280119７75.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级甘肃省一万名考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=280119７75. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年甘肃省一万名考试 考式 答案=280119７75.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级甘肃省一万名考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=280119７75人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”280119７75.祈福2015年甘肃省一万名考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级甘肃省一万名考试/ J7 J' y9 ]5 c5 w; D答案=280119７75.祈福2015年甘肃省一万名考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级甘肃省一万名考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年甘肃省一万名考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案280119７75.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=280119７75人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年甘肃省一万名考试 答案Ｑ280119７75"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15326293&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-07-10
其他媒体|1897620604|hefei|合肥专区|ZHO|2015-07-10 00:55:01|2015年河南特岗教师考试题 答案《★280119７75★》考后付|"2015年河南特岗教师考试题 答案《★280119７75★》考后付  2015年河南特岗教师考试 答案【通过率100%卡卡客服Ｑ280119７75包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年河南特岗教师考试真题答案-2015年河南特岗教师试题及 答案-2015年河南特岗教师考试时间-2015年河南特岗教师进村进社考试科目-2015年河南特岗教师考试大纲-2015年河南特岗教师考前答案-2015年河南特岗教师答案【Q280119７75包过】-2015年甘肃省一万名考试资料【Q280119７75包过】-2015年河南特岗教师复习资料-2015年河南特岗教师考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级河南特岗教师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年河南特岗教师考试 答案=280119７75- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级河南特岗教师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年河南特岗教师考试 答案 试题 真题 时间 科目〃Ｑ280119７75 ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年河南特岗教师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年甘肃省一万名考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案280119７75.祈福2015年内蒙古会计从业资ac格考试 考式 答案=280119７75+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级河南特岗教师考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=280119７75人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级河南特岗教师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级河南特岗教师考试 答案=280119７75.祈福2015年河南特岗教师进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年河南特岗教师考试 考式 答案=280119７75.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年河南特岗教师考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=280119７75人时简累 会受苦 正高级高级河南特岗教师考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=280119７75.祈福2015年河南特岗教师考试 考式 答案=280119７75人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级河南特岗教师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=280119７75.祈福2015年甘肃省一万名考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=280119７75 ^1 q) ~# t: {/ h/ J【=280119７75.祈福2015年河南特岗教师考试 考式 答案=280119７75 W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年河南特岗教师考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. 280119７75[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年河南特岗教师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=280119７75.祈福2015年甘肃省一万名考试 考式 答案=280119７75人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级河南特岗教师考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=280119７75_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级河南特岗教师答案【Q280119７75】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级河南特岗教师考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=280119７75 2015年河南特岗教师考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年河南特岗教师考试 考式 答案=280119７75.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年河南特岗教师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=280119７75 2015年河南特岗教师考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级河南特岗教师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W280119７75=280119７75 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^280119７75_100%】哪个2015年河南特岗教师考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=280119７75人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年甘肃省一万名考试 考式 答案=280119７75.+ F; ~ C( X7 G$ ?$ I祈福2015年河南特岗教师考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年河南特岗教师考试 考式 答案=280119７75.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级河南特岗教师答案【Q280119７75】9 I' [+ v* p3 m' Q=280119７75⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级甘肃省一万名 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年河南特岗教师考试 考式 答案=280119７75.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级河南特岗教师考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=280119７75. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年河南特岗教师考试 考式 答案=280119７75.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级河南特岗教师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=280119７75人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”280119７75.祈福2015年河南特岗教师考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级河南特岗教师考试/ J7 J' y9 ]5 c5 w; D答案=280119７75.祈福2015年甘肃省一万名考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级河南特岗教师考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年河南特岗教师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案280119７75.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=280119７75人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年河南特岗教师考试 答案Ｑ280119７75"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15326351&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-07-10
其他媒体|1897636828|hefei|合肥专区|ZHO|2015-07-10 01:08:01|2015年黑龙江特岗教师考试题 答案《★280119７75★》考后付|"2015年黑龙江特岗教师考试题 答案《★280119７75★》考后付  2015年黑龙江特岗教师考试 答案【通过率100%卡卡客服Ｑ280119７75包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年黑龙江特岗教师考试真题答案-2015年黑龙江特岗教师试题及 答案-2015年黑龙江特岗教师考试时间-2015年黑龙江特岗教师进村进社考试科目-2015年黑龙江特岗教师考试大纲-2015年黑龙江特岗教师考前答案-2015年黑龙江特岗教师答案【Q280119７75包过】-2015年黑龙江特岗教师考试资料【Q280119７75包过】-2015年黑龙江特岗教师复习资料-2015年黑龙江特岗教师考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级黑龙江特岗教师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年黑龙江特岗教师考试 答案=280119７75- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级黑龙江特岗教师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年黑龙江特岗教师考试 答案 试题 真题 时间 科目〃Ｑ280119７75 ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年黑龙江特岗教师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年黑龙江特岗教师考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案280119７75.祈福2015年内蒙古会计从业资ac格考试 考式 答案=280119７75+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级黑龙江特岗教师考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=280119７75人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级黑龙江特岗教师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级黑龙江特岗教师考试 答案=280119７75.祈福2015年黑龙江特岗教师进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年黑龙江特岗教师考试 考式 答案=280119７75.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年黑龙江特岗教师考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=280119７75人时简累 会受苦 正高级高级黑龙江特岗教师考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=280119７75.祈福2015年黑龙江特岗教师考试 考式 答案=280119７75人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级黑龙江特岗教师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=280119７75.祈福2015年黑龙江特岗教师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=280119７75 ^1 q) ~# t: {/ h/ J【=280119７75.祈福2015年黑龙江特岗教师考试 考式 答案=280119７75 W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年黑龙江特岗教师考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. 280119７75[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年黑龙江特岗教师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=280119７75.祈福2015年黑龙江特岗教师考试 考式 答案=280119７75人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级黑龙江特岗教师考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=280119７75_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级黑龙江特岗教师答案【Q280119７75】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级黑龙江特岗教师考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=280119７75 2015年黑龙江特岗教师考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年黑龙江特岗教师考试 考式 答案=280119７75.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年黑龙江特岗教师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=280119７75 2015年黑龙江特岗教师考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级黑龙江特岗教师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W280119７75=280119７75 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^280119７75_100%】哪个2015年黑龙江特岗教师考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=280119７75人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年黑龙江特岗教师考试 考式 答案=280119７75.+ F; ~ C( X7 G$ ?$ I祈福2015年黑龙江特岗教师考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年黑龙江特岗教师考试 考式 答案=280119７75.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级黑龙江特岗教师答案【Q280119７75】9 I' [+ v* p3 m' Q=280119７75⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级黑龙江特岗教师 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年黑龙江特岗教师考试 考式 答案=280119７75.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级黑龙江特岗教师考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=280119７75. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年黑龙江特岗教师考试 考式 答案=280119７75.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级黑龙江特岗教师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=280119７75人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”280119７75.祈福2015年黑龙江特岗教师考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级黑龙江特岗教师考试/ J7 J' y9 ]5 c5 w; D答案=280119７75.祈福2015年黑龙江特岗教师考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级黑龙江特岗教师考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年黑龙江特岗教师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案280119７75.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=280119７75人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年黑龙江特岗教师考试 答案Ｑ280119７75"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15326361&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-07-10
其他媒体|1898152586|hefei|合肥专区|ZHO|2015-07-10 10:46:01|2015年甘肃一万名考试题 答案《★７********★》|"2015年甘肃一万名考试题 答案《★７********★》  2015年甘肃一万名考试 答案【通过率100%卡卡客服Ｑ７********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年甘肃一万名考试真题答案-2015年甘肃一万名试题及 答案-2015年甘肃一万名考试时间-2015年甘肃一万名进村进社考试科目-2015年甘肃一万名考试大纲-2015年甘肃一万名考前答案-2015年甘肃一万名答案【Q７********包过】-2015年甘肃一万名考试资料【Q７********包过】-2015年甘肃一万名复习资料-2015年甘肃一万名考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级甘肃一万名著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年甘肃一万名考试 答案=７********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级甘肃一万名考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年甘肃一万名考试 答案 试题 真题 时间 科目〃Ｑ７******** ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年甘肃一万名考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年甘肃一万名考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案７********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=７********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级甘肃一万名考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=７********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级甘肃一万名考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级甘肃一万名考试 答案=７********.祈福2015年甘肃一万名进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年甘肃一万名考试 考式 答案=７********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年甘肃一万名考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=７********人时简累 会受苦 正高级高级甘肃一万名考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=７********.祈福2015年甘肃一万名考试 考式 答案=７********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级甘肃一万名考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=７********.祈福2015年甘肃一万名考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=７******** ^1 q) ~# t: {/ h/ J【=７********.祈福2015年甘肃一万名考试 考式 答案=７******** W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年甘肃一万名考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. ７********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年甘肃一万名考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=７********.祈福2015年甘肃一万名考试 考式 答案=７********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级甘肃一万名考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=７********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级甘肃一万名答案【Q７********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级甘肃一万名考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=７******** 2015年甘肃一万名考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年甘肃一万名考试 考式 答案=７********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年甘肃一万名考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=７******** 2015年甘肃一万名考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级甘肃一万名考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W７********=７******** 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^７********_100%】哪个2015年甘肃一万名考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=７********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年甘肃一万名考试 考式 答案=７********.+ F; ~ C( X7 G$ ?$ I祈福2015年甘肃一万名考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年甘肃一万名考试 考式 答案=７********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级甘肃一万名答案【Q７********】9 I' [+ v* p3 m' Q=７********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级甘肃一万名 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年甘肃一万名考试 考式 答案=７********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级甘肃一万名考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=７********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年甘肃一万名考试 考式 答案=７********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级甘肃一万名考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=７********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”７********.祈福2015年甘肃一万名考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级甘肃一万名考试/ J7 J' y9 ]5 c5 w; D答案=７********.祈福2015年甘肃一万名考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级甘肃一万名考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年甘肃一万名考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案７********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=７********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年甘肃一万名考试 答案Ｑ７********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15326626&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-07-10
其他媒体|1898345303|hefei|合肥专区|ZHO|2015-07-10 12:46:01|2015年甘肃省10000名考试题 答案《★７********★》|"2015年甘肃省10000名考试题 答案《★７********★》  2015年甘肃省10000名考试 答案【通过率100%卡卡客服Ｑ７********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年甘肃省10000名考试真题答案-2015年甘肃省10000名试题及 答案-2015年甘肃省10000名考试时间-2015年甘肃省10000名进村进社考试科目-2015年甘肃省10000名考试大纲-2015年河北特岗教师招聘考前答案-2015年甘肃省10000名答案【Q７********包过】-2015年河北特岗教师招聘考试资料【Q７********包过】-2015年甘肃省10000名复习资料-2015年甘肃省10000名考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级甘肃省10000名著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年河北特岗教师招聘考试 答案=７********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级甘肃省10000名考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年甘肃省10000名考试 答案 试题 真题 时间 科目〃Ｑ７******** ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年甘肃省10000名考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年河北特岗教师招聘考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案７********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=７********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级甘肃省10000名考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=７********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级河北特岗教师招聘考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级甘肃省10000名考试 答案=７********.祈福2015年甘肃省10000名进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年甘肃省10000名考试 考式 答案=７********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年河北特岗教师招聘考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=７********人时简累 会受苦 正高级高级甘肃省10000名考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=７********.祈福2015年甘肃省10000名考试 考式 答案=７********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级甘肃省10000名考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=７********.祈福2015年河北特岗教师招聘考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=７******** ^1 q) ~# t: {/ h/ J【=７********.祈福2015年甘肃省10000名考试 考式 答案=７******** W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年甘肃省10000名考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. ７********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年甘肃省10000名考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=７********.祈福2015年河北特岗教师招聘考试 考式 答案=７********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级河北特岗教师招聘考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=７********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级甘肃省10000名答案【Q７********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级甘肃省10000名考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=７******** 2015年甘肃省10000名考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年甘肃省10000名考试 考式 答案=７********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年甘肃省10000名考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=７******** 2015年甘肃省10000名考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级甘肃省10000名考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W７********=７******** 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^７********_100%】哪个2015年甘肃省10000名考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=７********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年河北特岗教师招聘考试 考式 答案=７********.+ F; ~ C( X7 G$ ?$ I祈福2015年甘肃省10000名考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年甘肃省10000名考试 考式 答案=７********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级甘肃省10000名答案【Q７********】9 I' [+ v* p3 m' Q=７********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级河北特岗教师招聘 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年甘肃省10000名考试 考式 答案=７********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级甘肃省10000名考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=７********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年甘肃省10000名考试 考式 答案=７********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级甘肃省10000名考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=７********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”７********.祈福2015年甘肃省10000名考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级甘肃省10000名考试/ J7 J' y9 ]5 c5 w; D答案=７********.祈福2015年河北特岗教师招聘考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级甘肃省10000名考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年甘肃省10000名考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案７********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=７********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年甘肃省10000名考试 答案Ｑ７********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15327106&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-07-10
其他媒体|1924650157|zhidao_baidu|电脑/网络 > 笔记本电脑|ZHO|2015-07-25 22:42:01|macbook pro 2015 13寸和 外星人 15最低配选哪个？？|macbook pro 2015 13寸和 外星人 15最低配选哪个？？4 分钟前格兰德法泽尓分类：苹果笔记本悬赏：10Mac戴尔笔记本笔记本电脑美留求问选哪现问题四：1、外星便携性底我知道3kg毕竟没手2、mbp装win底游戏性差要装win机器发热能否玩型游戏2k3、两种电脑性价比都低底哪款更低点4、两款质量问题断求神给高建|http://zhidao.baidu.com/question/1575624583932978820.html?entry=qb_browse_default|2015-07-25
其他媒体|1960159165|difang CN|地方频道 > 滚动读报|ZHO|2015-08-15 15:18:01|车界小鲜肉　k3s型动无极限|"最近|小鲜肉宁泽涛|于世锦赛男子100米自由泳决赛一举夺冠|向世界展示出“中国ing”的运动奇迹|赢得一片喝彩。明明可以靠颜值|却偏要拼实力的案例不止发生于体育赛场。在车市|秉承东风悦达起亚优质造车理念的k3s|拥有型格出众的外形设计和性能越级的巅峰实力|以“型动随我”的产品内涵|同样挑战着五门掀背车型的传统格局。作为东风悦达起亚旗下的风尚标杆|k3s以“简约直线美学”为设计理念|整体形象时尚动感。k3s有着张扬的宽大进气口|前中网则狭长精致|两者相辅相成；从侧面看|一条流畅的腰线贯穿首尾|传递出k3s极强的力量感；尾灯造型立体、饱满|极具辨识度的led后尾灯组合和镀铬饰条|锻造出豪华的品质感和高贵感。本稿件所含文字、图片和音视频资料 版权均属齐鲁晚报所有 任何媒体、网站或个人未经授权不得转载 违者将依法追究责任。"|http://difang.gmw.cn/newspaper/2015-08/15/content_108598583.htm|2015-08-15
其他媒体|1960237499|zhidao_baidu|生活 > 生活常识|ZHO|2015-08-15 16:29:01|东风悦达起亚k3保险杠4s店换还须要喷一到漆我|来自：手机知道汽车东风悦达起亚k3保险杠4s店换还须要喷一到漆我|http://zhidao.baidu.com/question/305544537022920564.html?fr=qlquick&entry=qb_list_default|2015-08-15
其他媒体|1970306917|difang CN|地方频道 > 滚动读报|ZHO|2015-08-21 09:06:01|ctcc南征肇庆 k3s技压群雄|烽火重燃 狼烟再起。8月16日 ctcc中国房车锦标赛第五站重回广东肇庆。在超级量产车组的冠军争夺战中 经过21圈的鏖战 东风悦达起亚车队小将张志强在最后一圈逆转取胜 携k3s赛车第二个冲过终点 跃居车手积分榜榜首 并帮助东风悦达起亚车队再次收获厂商杯冠军 继续领跑超级量产车组。在ctcc已完成的五站比赛中 东风悦达起亚车队曾多次上演绝地反击 除了车手的出色发挥 k3s赛车的优异品质亦功不可没。一个汽车品牌的荣耀 在于赢得赛场的同时 更能赢得消费者的坚定追随。承袭东风悦达起亚k系家族血脉的k3s 必将持续创造市场与赛道荣誉的双丰收。|http://difang.gmw.cn/newspaper/2015-08/21/content_108723173.htm|2015-08-21
其他媒体|1978565959|difang CN|地方频道 > 滚动读报|ZHO|2015-08-26 03:53:01|k3s征战ctcc再夺冠|8月16日 ctcc中国房车锦标赛第五站重回广东肇庆。在超级量产车组的冠军争夺战中 经过21圈的鏖战 东风悦达起亚车队小将张志强在最后一圈逆转取胜 携k3s赛车第二个冲过终点 跃居车手积分榜榜首 并帮助东风悦达起亚车队再次收获厂商杯冠军 继续领跑超级量产车组。在ctcc已完成的五站比赛中 东风悦达起亚车队曾多次上演绝地反击 除了车手的出色发挥之外 k3s赛车的品质也功不可没。其搭载的1.6t-gdi发动机 是由1.6tgdigamma发动机升级改装而来 并因ctcc赛场需求进一步升级 达到了310马力。此外 k3s赛车的操控性和稳定性不仅“擅长”直线加速 更有精彩的弯道表现。值得一提的是 k3s赛车发动机是由起亚技术中心自主研发 彰显出东风悦达起亚在另一条“技术战线”上 同样具备强大的竞争优势。(黄天姣）|http://difang.gmw.cn/newspaper/2015-08/26/content_108812286.htm|2015-08-26
其他媒体|1978621661|difang CN|地方频道 > 滚动读报|ZHO|2015-08-26 05:23:02|一卡玩转三镇健身场馆|本报记者李勇为推进全民健身运动 为实现都市圈“健身一卡通”计划 长江日报报业集团下属子媒《武汉商报》联合光大银行于6月18日正式启动“大武汉健身联盟” 只需499元/年 即可在二十余家跨区健身会所健身 还有“299元季卡” 可通用十余家游泳及羽毛球馆。自从消息见报后 吸引了众多市民的关注 健身爱好者、公司员工、大学毕业生 纷纷拨打咨询电话详细询问后 立刻加入这一联盟 玩转三镇的健身场馆。今年大学刚刚毕业的晶晶这个暑假过得不一般 没有像师哥师姐那样在炎炎夏日下 四处奔波辛苦地找工作 晶晶给自己制定了一个计划 一边找工作一边健身锻炼。在得知有“大武汉健身联盟”后 晶晶和同学不久前一起到附近的光大银行营业点 很方便的就办理一张大武汉健身联盟卡。平时 她们总是把卡随身携带 在汉口面试完了 就在汉口的健身房练练瑜伽 放松放松心情；在武昌面试完了后 就在武昌找家游泳馆学习游泳；在汉阳面试完了后 就在汉阳打一场愉快的羽毛球。辛苦而紧张的面试历程 在晶晶和同学的眼里变得既轻松又愉快。在接受采访时 她笑着表示 有了健康完美的身体 自然好找工作哦。大武汉健身联盟场馆序号场馆名称地址类别1艾思特健身中心(st健身)武昌区彭刘杨西路汉飞逛逛街1号楼4楼(武汉音乐学院)年卡2菲力健身俱乐部汉口大智路轻轨站黄兴路沃尔玛二楼年卡3飞运动国际健身俱乐部（南湖店）武昌凯旋名邸商铺年卡4武汉市武昌区新韵动健身工作室洪山区徐东大街120号福星惠誉群星城k3-2702室年卡5格美健身俱乐部（后湖店）江岸区后湖二路与兴业南路交界口（中百超市二楼）年卡6帝斯力高级私人健身会所武昌中北路124号德成中心27楼年卡7彩虹健身（原超级健身）花桥街天成花园1号楼1栋2楼（豪泰宾馆二楼）年卡8斯巴达健身私教会所汉阳区汉阳大道闽东国际商业西区3楼2室（家乐福旁）年卡9三角湖羽毛球馆汉阳东风大道83号（经开万达对面）年卡10道义（嘉禾园）健身俱乐部东西湖区一清路嘉禾园小区内年卡11琥珀健身馆武昌区积玉桥万达soho12号楼3楼季卡12水立方游泳馆水立方商务会馆后湖大道99号季卡13保利大酒店游泳馆武昌区民主路788号季卡14天天游泳馆汉阳区芳草路88号（龙阳1号内）季卡15月亮湾游泳馆武昌区临江大道三层楼站(武昌热电厂对面)季卡16七一游泳馆京汉大道七一中学旁季卡17长城羽毛球馆江汉区建设大道575号（贵宾楼与加油站中间进去100米）季卡18英弢羽毛球馆京汉大道259号附近季卡19百利羽毛球馆武昌区徐东大街88号麦德龙后面季卡20翔云羽毛球馆江岸区解放大道2020号（丹水池天桥旁中国储运院内）季卡21天天羽毛球馆汉阳区龙阳大道康大路5号季卡22奥林乒乓球俱乐部江汉区振兴路72号季卡23羽乐羽毛球馆武昌洪山区图书城18号（瑞安王朝酒店附近）季卡办卡方式报名热线：027-*******、027-*******报名地址：长江日报路2号（长江日报内）、武汉市内光大银行各营业网点加盟电话：*******（孙）上周读者报名踊跃 200份礼品已经送完 现为满足广大读者的要求 增加200个名额。即日起 办理499元年卡 前200名报名读者送：●价值299元季卡●价值888元兰丁（国际）健康体检管理中心提供的专业体检套餐1次●价值150元“一号蓝”有机野生草莓汁一箱|http://difang.gmw.cn/newspaper/2015-08/26/content_108813707.htm|2015-08-26
其他媒体|1978817096|zhidao_baidu|电脑/网络 > 硬件 > 硬盘|ZHO|2015-08-26 09:28:01|请问广汽本田锋范手动精英版跟东风悦达k3谁比较好点|来自：手机知道汽车|http://zhidao.baidu.com/question/1176840476375317259.html?fr=qlquick&entry=qb_list_default|2015-08-26
其他媒体|1979257317|hefei|合肥专区|ZHO|2015-08-26 14:22:02|2015年安全工程师考试 答案《★*********★》|"2015年安全工程师考试 答案《★*********★》  2015年安全工程师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年安全工程师考试真题答案-2015年安全工程师试题及 答案-2015年安全工程师考试时间-2015年安全工程师进村进社考试科目-2015年安全工程师考试大纲-2015年安全工程师考前答案-2015年安全工程师答案【Q*********包过】-2015年安全工程师考试资料【Q*********包过】-2015年安全工程师复习资料-2015年安全工程师考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级安全工程师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年安全工程师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级安全工程师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年安全工程师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年安全工程师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年安全工程师考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级安全工程师考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级安全工程师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级安全工程师考试 答案=*********.祈福2015年安全工程师进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年安全工程师考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年安全工程师考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级安全工程师考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年安全工程师考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级安全工程师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年安全工程师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年安全工程师考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年安全工程师考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年安全工程师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年安全工程师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级安全工程师考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级安全工程师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级安全工程师考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年安全工程师考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年安全工程师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年安全工程师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年安全工程师考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级安全工程师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年安全工程师考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年安全工程师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年安全工程师考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年安全工程师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级安全工程师答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级安全工程师 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年安全工程师考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级安全工程师考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年安全工程师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级安全工程师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年安全工程师考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级安全工程师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年安全工程师考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级安全工程师考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年安全工程师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年安全工程师考试 答案Ｑ*********2015年安全工程师考试 答案《★*********★》"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15494682&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-08-26
其他媒体|1979257320|hefei|合肥专区|ZHO|2015-08-26 14:22:03|2015年暖通工程师考试 答案《★*********★》|"2015年暖通工程师考试 答案《★*********★》  2015年暖通工程师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年暖通工程师考试真题答案-2015年暖通工程师试题及 答案-2015年暖通工程师考试时间-2015年暖通工程师进村进社考试科目-2015年暖通工程师考试大纲-2015年暖通工程师考前答案-2015年暖通工程师答案【Q*********包过】-2015年暖通工程师考试资料【Q*********包过】-2015年暖通工程师复习资料-2015年暖通工程师考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级暖通工程师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年暖通工程师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级暖通工程师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年暖通工程师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年暖通工程师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年暖通工程师考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级暖通工程师考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级暖通工程师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级暖通工程师考试 答案=*********.祈福2015年暖通工程师进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年暖通工程师考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年暖通工程师考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级暖通工程师考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年暖通工程师考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级暖通工程师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年暖通工程师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年暖通工程师考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年暖通工程师考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年暖通工程师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年暖通工程师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级暖通工程师考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级暖通工程师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级暖通工程师考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年暖通工程师考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年暖通工程师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年暖通工程师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年暖通工程师考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级暖通工程师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年暖通工程师考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年暖通工程师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年暖通工程师考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年暖通工程师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级暖通工程师答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级暖通工程师 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年暖通工程师考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级暖通工程师考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年暖通工程师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级暖通工程师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年暖通工程师考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级暖通工程师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年暖通工程师考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级暖通工程师考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年暖通工程师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年暖通工程师考试 答案Ｑ*********2015年暖通工程师考试 答案《★*********★》"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15494899&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-08-26
其他媒体|1979297054|hefei|合肥专区|ZHO|2015-08-26 14:48:01|2015年注安考试 答案《★*********★》|"2015年注安考试 答案《★*********★》  2015年注安考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年注安考试真题答案-2015年注安试题及 答案-2015年注安考试时间-2015年注安进村进社考试科目-2015年注安考试大纲-2015年注安考前答案-2015年注安答案【Q*********包过】-2015年注安考试资料【Q*********包过】-2015年注安复习资料-2015年注安考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级注安著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年注安考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级注安考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年注安考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年注安考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年注安考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级注安考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级注安考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级注安考试 答案=*********.祈福2015年注安进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年注安考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年注安考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级注安考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年注安考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级注安考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年注安考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年注安考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年注安考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年注安考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年注安考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级注安考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级注安答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级注安考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年注安考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年注安考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年注安考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年注安考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级注安考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年注安考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年注安考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年注安考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年注安考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级注安答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级注安 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年注安考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级注安考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年注安考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级注安考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年注安考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级注安考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年注安考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级注安考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年注安考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年注安考试 答案Ｑ*********2015年注安考试 答案《★*********★》"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15494426&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-08-26
其他媒体|1979297055|hefei|合肥专区|ZHO|2015-08-26 14:48:01|2015年给排水工程师考试 答案《★*********★》|"2015年给排水工程师考试 答案《★*********★》  2015年给排水工程师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年给排水工程师考试真题答案-2015年给排水工程师试题及 答案-2015年给排水工程师考试时间-2015年给排水工程师进村进社考试科目-2015年给排水工程师考试大纲-2015年给排水工程师考前答案-2015年给排水工程师答案【Q*********包过】-2015年给排水工程师考试资料【Q*********包过】-2015年给排水工程师复习资料-2015年给排水工程师考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级给排水工程师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年给排水工程师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级给排水工程师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年给排水工程师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年给排水工程师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年给排水工程师考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级给排水工程师考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级给排水工程师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级给排水工程师考试 答案=*********.祈福2015年给排水工程师进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年给排水工程师考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年给排水工程师考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级给排水工程师考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年给排水工程师考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级给排水工程师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年给排水工程师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年给排水工程师考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年给排水工程师考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年给排水工程师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年给排水工程师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级给排水工程师考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级给排水工程师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级给排水工程师考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年给排水工程师考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年给排水工程师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年给排水工程师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年给排水工程师考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级给排水工程师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年给排水工程师考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年给排水工程师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年给排水工程师考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年给排水工程师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级给排水工程师答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级给排水工程师 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年给排水工程师考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级给排水工程师考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年给排水工程师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级给排水工程师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年给排水工程师考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级给排水工程师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年给排水工程师考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级给排水工程师考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年给排水工程师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年给排水工程师考试 答案Ｑ*********2015年给排水工程师考试 答案《★*********★》"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15495137&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-08-26
其他媒体|1979297056|hefei|合肥专区|ZHO|2015-08-26 14:48:01|2015年电气工程师考试 答案《★*********★》|"2015年电气工程师考试 答案《★*********★》  2015年电气工程师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年电气工程师考试真题答案-2015年电气工程师试题及 答案-2015年电气工程师考试时间-2015年电气工程师进村进社考试科目-2015年电气工程师考试大纲-2015年电气工程师考前答案-2015年电气工程师答案【Q*********包过】-2015年电气工程师考试资料【Q*********包过】-2015年电气工程师复习资料-2015年电气工程师考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级电气工程师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年电气工程师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级电气工程师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年电气工程师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年电气工程师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年电气工程师考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级电气工程师考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级电气工程师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级电气工程师考试 答案=*********.祈福2015年电气工程师进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年电气工程师考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年电气工程师考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级电气工程师考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年电气工程师考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级电气工程师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年电气工程师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年电气工程师考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年电气工程师考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年电气工程师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年电气工程师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级电气工程师考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级电气工程师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级电气工程师考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年电气工程师考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年电气工程师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年电气工程师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年电气工程师考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级电气工程师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年电气工程师考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年电气工程师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年电气工程师考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年电气工程师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级电气工程师答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级电气工程师 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年电气工程师考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级电气工程师考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年电气工程师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级电气工程师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年电气工程师考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级电气工程师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年电气工程师考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级电气工程师考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年电气工程师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年电气工程师考试 答案Ｑ*********2015年电气工程师考试 答案《★*********★》"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15495247&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-08-26
其他媒体|1979297057|hefei|合肥专区|ZHO|2015-08-26 14:48:01|2015年岩土工程师考试 答案《★*********★》|"2015年岩土工程师考试 答案《★*********★》  2015年岩土工程师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年岩土工程师考试真题答案-2015年岩土工程师试题及 答案-2015年岩土工程师考试时间-2015年岩土工程师进村进社考试科目-2015年岩土工程师考试大纲-2015年岩土工程师考前答案-2015年岩土工程师答案【Q*********包过】-2015年岩土工程师考试资料【Q*********包过】-2015年岩土工程师复习资料-2015年岩土工程师考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级岩土工程师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年岩土工程师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级岩土工程师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年岩土工程师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年岩土工程师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年岩土工程师考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级岩土工程师考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级岩土工程师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级岩土工程师考试 答案=*********.祈福2015年岩土工程师进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年岩土工程师考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年岩土工程师考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级岩土工程师考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年岩土工程师考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级岩土工程师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年岩土工程师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年岩土工程师考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年岩土工程师考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年岩土工程师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年岩土工程师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级岩土工程师考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级岩土工程师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级岩土工程师考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年岩土工程师考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年岩土工程师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年岩土工程师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年岩土工程师考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级岩土工程师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年岩土工程师考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年岩土工程师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年岩土工程师考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年岩土工程师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级岩土工程师答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级岩土工程师 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年岩土工程师考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级岩土工程师考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年岩土工程师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级岩土工程师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年岩土工程师考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级岩土工程师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年岩土工程师考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级岩土工程师考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年岩土工程师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年岩土工程师考试 答案Ｑ*********2015年岩土工程师考试 答案《★*********★》"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15495264&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-08-26
其他媒体|1979297058|hefei|合肥专区|ZHO|2015-08-26 14:48:01|2015年化工工程师考试 答案《★*********★》|"2015年化工工程师考试 答案《★*********★》  2015年化工工程师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年化工工程师考试真题答案-2015年化工工程师试题及 答案-2015年化工工程师考试时间-2015年化工工程师进村进社考试科目-2015年化工工程师考试大纲-2015年化工工程师考前答案-2015年化工工程师答案【Q*********包过】-2015年化工工程师考试资料【Q*********包过】-2015年化工工程师复习资料-2015年化工工程师考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级化工工程师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年化工工程师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级化工工程师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年化工工程师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年化工工程师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年化工工程师考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级化工工程师考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级化工工程师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级化工工程师考试 答案=*********.祈福2015年化工工程师进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年化工工程师考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年化工工程师考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级化工工程师考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年化工工程师考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级化工工程师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年化工工程师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年化工工程师考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年化工工程师考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年化工工程师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年化工工程师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级化工工程师考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级化工工程师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级化工工程师考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年化工工程师考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年化工工程师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年化工工程师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年化工工程师考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级化工工程师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年化工工程师考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年化工工程师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年化工工程师考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年化工工程师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级化工工程师答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级化工工程师 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年化工工程师考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级化工工程师考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年化工工程师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级化工工程师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年化工工程师考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级化工工程师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年化工工程师考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级化工工程师考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年化工工程师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年化工工程师考试 答案Ｑ*********2015年化工工程师考试 答案《★*********★》"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15495279&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-08-26
其他媒体|1979297059|hefei|合肥专区|ZHO|2015-08-26 14:48:01|2015年环保工程师考试 答案《★*********★》|"2015年环保工程师考试 答案《★*********★》  2015年环保工程师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年环保工程师考试真题答案-2015年环保工程师试题及 答案-2015年环保工程师考试时间-2015年环保工程师进村进社考试科目-2015年环保工程师考试大纲-2015年环保工程师考前答案-2015年环保工程师答案【Q*********包过】-2015年环保工程师考试资料【Q*********包过】-2015年环保工程师复习资料-2015年环保工程师考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级环保工程师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年环保工程师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级环保工程师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年环保工程师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年环保工程师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年环保工程师考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级环保工程师考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级环保工程师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级环保工程师考试 答案=*********.祈福2015年环保工程师进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年环保工程师考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年环保工程师考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级环保工程师考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年环保工程师考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级环保工程师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年环保工程师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年环保工程师考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年环保工程师考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年环保工程师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年环保工程师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级环保工程师考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级环保工程师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级环保工程师考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年环保工程师考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年环保工程师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年环保工程师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年环保工程师考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级环保工程师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年环保工程师考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年环保工程师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年环保工程师考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年环保工程师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级环保工程师答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级环保工程师 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年环保工程师考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级环保工程师考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年环保工程师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级环保工程师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年环保工程师考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级环保工程师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年环保工程师考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级环保工程师考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年环保工程师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年环保工程师考试 答案Ｑ*********2015年环保工程师考试 答案《★*********★》"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15495304&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-08-26
其他媒体|1979297060|hefei|合肥专区|ZHO|2015-08-26 14:48:01|2015年一级结构工程师考试 答案《★*********★》|"2015年一级结构工程师考试 答案《★*********★》  2015年一级结构工程师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年一级结构工程师考试真题答案-2015年一级结构工程师试题及 答案-2015年一级结构工程师考试时间-2015年一级结构工程师进村进社考试科目-2015年一级结构工程师考试大纲-2015年一级结构工程师考前答案-2015年一级结构工程师答案【Q*********包过】-2015年一级结构工程师考试资料【Q*********包过】-2015年一级结构工程师复习资料-2015年一级结构工程师考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级一级结构工程师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年一级结构工程师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级一级结构工程师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年一级结构工程师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年一级结构工程师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年一级结构工程师考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级一级结构工程师考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级一级结构工程师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级一级结构工程师考试 答案=*********.祈福2015年一级结构工程师进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年一级结构工程师考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年一级结构工程师考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级一级结构工程师考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年一级结构工程师考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级一级结构工程师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年一级结构工程师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年一级结构工程师考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年一级结构工程师考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年一级结构工程师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年一级结构工程师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级一级结构工程师考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级一级结构工程师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级一级结构工程师考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年一级结构工程师考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年一级结构工程师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年一级结构工程师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年一级结构工程师考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级一级结构工程师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年一级结构工程师考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年一级结构工程师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年一级结构工程师考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年一级结构工程师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级一级结构工程师答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级一级结构工程师 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年一级结构工程师考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级一级结构工程师考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年一级结构工程师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级一级结构工程师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年一级结构工程师考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级一级结构工程师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年一级结构工程师考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级一级结构工程师考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年一级结构工程师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年一级结构工程师考试 答案Ｑ*********2015年一级结构工程师考试 答案《★*********★》"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15495324&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-08-26
其他媒体|1979297061|hefei|合肥专区|ZHO|2015-08-26 14:48:01|2015年价格鉴证师考试 答案《★*********★》|"2015年价格鉴证师考试 答案《★*********★》  2015年价格鉴证师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年价格鉴证师考试真题答案-2015年价格鉴证师试题及 答案-2015年价格鉴证师考试时间-2015年价格鉴证师进村进社考试科目-2015年价格鉴证师考试大纲-2015年价格鉴证师考前答案-2015年价格鉴证师答案【Q*********包过】-2015年价格鉴证师考试资料【Q*********包过】-2015年价格鉴证师复习资料-2015年价格鉴证师考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级价格鉴证师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年价格鉴证师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级价格鉴证师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年价格鉴证师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年价格鉴证师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年价格鉴证师考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级价格鉴证师考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级价格鉴证师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级价格鉴证师考试 答案=*********.祈福2015年价格鉴证师进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年价格鉴证师考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年价格鉴证师考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级价格鉴证师考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年价格鉴证师考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级价格鉴证师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年价格鉴证师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年价格鉴证师考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年价格鉴证师考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年价格鉴证师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年价格鉴证师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级价格鉴证师考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级价格鉴证师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级价格鉴证师考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年价格鉴证师考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年价格鉴证师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年价格鉴证师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年价格鉴证师考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级价格鉴证师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年价格鉴证师考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年价格鉴证师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年价格鉴证师考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年价格鉴证师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级价格鉴证师答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级价格鉴证师 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年价格鉴证师考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级价格鉴证师考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年价格鉴证师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级价格鉴证师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年价格鉴证师考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级价格鉴证师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年价格鉴证师考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级价格鉴证师考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年价格鉴证师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年价格鉴证师考试 答案Ｑ*********2015年价格鉴证师考试 答案《★*********★》"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15495408&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-08-26
其他媒体|1979297062|hefei|合肥专区|ZHO|2015-08-26 14:48:01|2015年二级结构工程师考试 答案《★*********★》|"2015年二级结构工程师考试 答案《★*********★》  2015年二级结构工程师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年二级结构工程师考试真题答案-2015年二级结构工程师试题及 答案-2015年二级结构工程师考试时间-2015年二级结构工程师进村进社考试科目-2015年二级结构工程师考试大纲-2015年二级结构工程师考前答案-2015年二级结构工程师答案【Q*********包过】-2015年二级结构工程师考试资料【Q*********包过】-2015年二级结构工程师复习资料-2015年二级结构工程师考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级二级结构工程师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年二级结构工程师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级二级结构工程师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年二级结构工程师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年二级结构工程师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年二级结构工程师考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级二级结构工程师考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级二级结构工程师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级二级结构工程师考试 答案=*********.祈福2015年二级结构工程师进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年二级结构工程师考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年二级结构工程师考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级二级结构工程师考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年二级结构工程师考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级二级结构工程师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年二级结构工程师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年二级结构工程师考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年二级结构工程师考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年二级结构工程师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年二级结构工程师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级二级结构工程师考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级二级结构工程师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级二级结构工程师考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年二级结构工程师考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年二级结构工程师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年二级结构工程师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年二级结构工程师考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级二级结构工程师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年二级结构工程师考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年二级结构工程师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年二级结构工程师考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年二级结构工程师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级二级结构工程师答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级二级结构工程师 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年二级结构工程师考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级二级结构工程师考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年二级结构工程师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级二级结构工程师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年二级结构工程师考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级二级结构工程师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年二级结构工程师考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级二级结构工程师考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年二级结构工程师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年二级结构工程师考试 答案Ｑ*********2015年二级结构工程师考试 答案《★*********★》"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15495457&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-08-26
其他社区|1980043864|yam|即時 > 宅趣|ZHO|2015-08-26 22:33:02|韓國CGV電影院可自製《照片票根》把票根用拍立得方式收藏起來♥|圖片來自：instagram.com/chan_hyeok316不少人都會收藏票根做紀念 尤其跟另一半出遊更喜歡把大小收據留著 做為當次約會的回憶。不過票券留久會開始泛黃 如果是熱感應紙收據還會因久放的關係讓上面文字消失 想拿出來回味才發現剩白紙一張T^T韓國連鎖電影院CGV就提供一項特別服務 可以把你的票根用照片方式印出變成照片票根 瞬間讓收藏值爆增！  在社群上只要搜尋포토티켓就有很多照片票根的美照 韓國民眾對於可以用照片方式保存票根表示非常滿意～(笑)  圖片來自：instagram.co... 【文章內容不代表蕃薯藤立場 想看更多歡迎到>>>卡卡洛普－宅宅新聞】     蕃Plus+1+1     -->|http://n.yam.com/gamme/otaku/20150826/20150826239534.html|2015-08-26
其他媒体|2039011239|zhidao_baidu|烦恼|ZHO|2015-10-01 00:26:03|东风悦达起亚k3一月销售多少辆|来自：手机知道汽车|http://zhidao.baidu.com/question/265344175614285485.html?fr=qlquick&entry=qb_list_default|2015-10-01
各大媒体|2039534197|chinanews|时政经济|ZHO|2015-10-01 10:07:03|陕西交警权威发布十一最全出行攻略|您的位置：首页   时政经济 	 陕西交警权威发布十一最全出行攻略    2015年10月01日 08:39   来源：   西部网    	               	 　　十一黄金周将至 受高速公路免费刺激 外出旅游和自驾游人群激增 道路交通压力剧增 针对陕西省内道路状况 省公安厅交警总队发布五大类交通出行提示 让市民提前获悉出行信息 避免不必要的拥堵。　　同时 交警部门提醒全省广大群众 出行前应该提前了解出行目的地的交通状况 做好安排。如果遇到拥堵和事故路段时请听从交警指挥 一旦车辆发生故障或事故 应保护好事故现场 及时拨打122报警 对于刮蹭等轻微事故则建议走快速理赔。　　一、陕西全省高速公路限速提示　　1、连霍高速陕西段(G30)：渭南潼关至宝鸡段 途经华阴、华县、渭南、西安、咸阳、兴平、武功、杨凌、扶风、眉县 限速110Km/h(双向四车道)-120Km/h(双向八车道) 宝鸡至陈仓省际站 最高限速80Km/h 其中隧道最高限速60Km/h。绕城高速阿房宫收费站至兴平段 限速120Km/h。　　2、包茂高速陕西段(G65)：西安至榆林段 途经高陵、三原、铜川、宜君、黄陵、洛川、富县、甘泉、延安、安塞、靖边、横山 限速80Km/h(山区段)-100Km/h(平川段) 西安至安康段 途经柞水、镇安、安康、紫阳 限速80Km/h(山区段)-100Km/h(平川段) 其中隧道最高限速60Km/h。　　延西高速(G65W)西安至铜川段 限速120 Km/h。　　3、福银高速陕西段(G70)：西长段 途经咸阳、礼泉、乾县、永寿、彬县、长武 限速80Km/h-120Km/h 西商、商漫段 途经蓝田、商洛、山阳 限速80Km/h-100Km/h其中隧道限速60Km/h。　　4、沪陕高速陕西段(G40)：西安至蓝田段 限速120Km/h；商洛段 途经商洛、丹凤、商南 限速80Km/h- 100Km/h 其中隧道最高限速60Km/h。　　5、京昆高速陕西段(G5)：西禹段 途经高陵、阎良、富平、澄城、合阳、韩城 限速120Km/h；西汉段 途户县、宁陕、佛坪、洋县 限速80Km/h(山区)-120Km/h 隧道最高限速60Km/h。汉宁段 途经洋县、城固、汉中、南郑、勉县、宁强 限速80Km/h-100Km/h 隧道最高限速60Km/h。　　6、青银高速陕西段(G20)：途经吴堡、绥德、子洲、横山、靖边、定边 限速80Km/h-100Km/h。　　7、青兰高速陕西段(G22)：途经壶口、宜川、富县 限速80Km/h-100Km/h 隧道最高限速60Km/h。　　8、十天高速陕西段(G7011)：途经白河、旬阳、安康、汉阴、石泉、西乡、汉中、勉县、略阳 限速80Km/h-100Km/h 隧道限速60 Km/h。　　二、陕西境内高速事故多发路段及安全提示　　1、京昆高速陕西段(G5)：渭南境内澄城韦庄段连续坡道加弯道；西安境内涝峪口至秦岭1号隧道段为山区高速 弯多、坡陡、桥隧相连 易发生追尾事故；汉中境内铁炉沟隧道内视线不良 弯道连续下坡。　　2、沪陕高速陕西段(G40)：西安境内蓝田段、商洛境内商南段山区高速 弯道多、纵坡大、桥隧相连。　　安全提醒：在上述路段行驶时 严格遵守限速标准 保持安全车距、平稳驾驶 避免长时间连续使用刹车。遇道路湿滑等情况 应平稳降低车速 握紧方向 避免急刹车、急打方向；进入隧道前要及时打开车灯 降低车速 注意观察 谨慎通过。　　3、316国道：安康旬阳境内吕河大桥北 该路段属于三级道路 路面较窄 紧邻汉江 易发生车辆翻坠或撞崖事故。　　安全提醒：驾车经过上述路段时 一定不要超速、超载行驶 还要避免超车、随意变道 切不可连续使用刹车 严禁占道停车 保持安全车距 依次通过。　　4、107省道：西安市长安区境内道路 沿途遍布村庄、旅游景点、农家乐 上百个平交道口与107省道相连。且沿途汽车、摩托车、低速载货汽车、拖拉机、非机动车、行人等混行 沿途摆摊设点较多 交通环境复杂 极易发生汽车碰撞摩托车、非机动车、行人的交通事故。　　安全提醒：驾车经过此路段时。要降低车速、减速慢行 经过平交道口要注意观察是否有行人通过 并鸣笛提示。　　三、全省高速公路施工情况　　1、西安绕城高速：杏园立交改扩建施工 道路通行阻塞(施工导致上、下行各两个车道通行)；尚航璐下穿绕城高速施工因后期路面恢复 暂时通行阻塞(单幅双向通行 各保证两个车道通行)。　　2、沪陕高速西商段：洛岔高速洛南方向下行k2+900米处护坡施工 k0+800米至k3+400米处实行单幅双向通行。因渭南至玉山高速公路施工需要 国庆期间西安方向上行k1478+600米至上行k1480+800米封闭第三车道、紧急停车带 一、二车道正常通行；商洛方向下行k1481+800米至下行k1480+100米封闭第三车道、紧急停车带 一、二车道正常通行。　　3、沪陕高速商界段：因比亚迪东西厂区修建连接通道 沪陕商洛东收费站出入口连接线k140至k180之间占道施工 请过往车辆按照交通指示绕行西侧便道通行。　　4、包茂高速安川段：包茂高速小康段下行k1074+100处郑家湾2#桥进行施工。施工期间在上行k1073+600米至上行k1074+200米出实施单幅双向通车的方式进行保畅 施工期间途经此路段车辆 请严格按照现场标识标线行驶。　　5、包茂高速延靖段：黄延高速公路(在建)k534+360---k536+830与包茂高速公路(延靖段)马家沟枢纽拼接路面施工 占用应急车道 严格要求施工单位按照《公路养护安全作业规程》摆放施工标志标牌 施工区增设围挡 陆正加强施工监管。　　6、青兰高速宜富段：2015年9月1日至2015年10月15日往雷家角方向直落隧道封闭施工 宜富高速k1224+500米至k1227+400米 实行单幅双向通行；2015年9月8 日至2015年10月15 日往壶口方向石家河隧道封闭施工 宜富高速k1187+700至k1190+500实行单幅双向通行；2015年9月12 日至2015年10月15日往壶口方向吉家村隧道封闭施工 宜富高速k1177+700至k1182+ooo实行单幅双向通行。　　7、延志吴高速：因进行隧道检测 延志吴高速志丹东隧道上行线延安至志丹方向全部封闭 志丹东隧道下行线志丹至延安方向k46+150m---k51+450m处实行单幅双向通行；马鞍子隧道下行线吴起至延安方向k106+756m---k106+786m处进行路基病害处理工程 占用行车道。　　8、榆神高速：榆神高速神木至店塔段k57+260处进行神木县第二新村至西过境路连接大桥上跨桥梁施工 施工期间实行单幅双向通行；双向禁止宽度超过5米的货车通行；请过往车辆严格按照施工指示标志 减速慢行。　　9、G30连霍高速西安至渭南段：因改扩建施工 连霍高速西临段全线禁止7座以上(不含7座)客车及货车通行 7座以下客车单幅双向通行；灞桥收费站入口禁止7座以上客车及货车通行 临潼、豁口收费站出入口禁止所有车辆通行。兵马俑专线将实施交通管制 禁止7座(不含7座)以上客车及货车驶入。前往兵马俑的7座以上客车及货车 可从兵马俑邻近的新丰收费站驶出高速 绕行G310国道到达。受西临高速施工影响西渭段新丰、兵马俑收费站入口往西安方向禁止7座以上客车及货车通行。　　四、旅游景区道路及安全提示　　1、秦始皇兵马俑博物馆：位于距西安27公里的临潼区。路线：G30连霍高速西安??秦俑旅游专线兵??马俑收费站 到达景区。G30单幅双向通行；低速：G108双向四车道；因改扩建施工 连霍高速西临段全线禁止7座以上(不含7座)客车及货车通行 7座以下客车单幅双向通行；灞桥收费站入口禁止7座以上客车及货车通行 临潼、豁口收费站出入口禁止所有车辆通行。兵马俑专线将实施交通管制 禁止7座(不含7座)以上客车及货车驶入。前往兵马俑的7座以上客车及货车 可从兵马俑邻近的新丰收费站驶出高速 绕行G310国道到达。　受西临高速施工影响西渭段新丰、兵马俑收费站入口往西安方向禁止7座以上客车及货车通行。 　　2、唐华清宫 位于距西安27公里的临潼区。路线：G30连霍高速西安??斜口收费站下高速??G108进入临潼城区至秦唐大道3km到达景区。低速：G108双向四车道进入临潼城区至秦唐大道3km到达景区。　　3、宝鸡法门寺 位于陕西省宝鸡市扶风县。距西安市110公里。距宝鸡市70公里。自驾游的旅客可通过G30(连霍高速)西安到宝鸡段通行。也可通行310国道或104省道到扶风县法门镇。另外 游客也可从西安市城西客运站乘坐长途客车前往。节日期间 无道路施工。路况良好。　　4、宝鸡太白山 位于陕西省宝鸡市眉县。距西安市110公里。距宝鸡市75公里。自驾游的旅客可通过G30(连霍高速)西安到宝鸡段通行。也可通行310国道到眉县汤浴镇。另外 游客也可从西安市乘坐长途客车前往。节日期间 无道路施工。路况良好。太白山景区禁止社会车辆通行。游客必须乘坐景区旅游车辆出入景区。　　5、宝鸡红河谷 位于陕西省宝鸡市眉县。距西安市120公里。距宝鸡市65公里。自驾游的旅客可通过G30(连霍高速)西安到宝鸡段通行。也可通行310国道到眉县金渠镇。另外 游客也可从西安市乘坐长途客车前往。节日期间 无道路施工。路况良好。　　6、宝鸡关山牧场 位于陕西省宝鸡市陇县。距西安市约300公里。距宝鸡市110公里。自驾游的旅客可通过G30(连霍高速)从西安到宝鸡 再转道宝平(宝鸡到平凉)高速通行。也可通行310国道到宝鸡后转道212省道或从西安通行104省道到陇县后转道景区专用线。另外 游客也可从西安市乘坐长途客车前往。节日期间 无道路施工。路况良好。关山牧场景区道路属于山区道路 弯道较多 请驾驶员朋友谨慎驾驶 切忌超速超员。　　7、咸阳马嵬驿 位于陕西省兴平市西约11公里。马嵬距西安咸阳机场约39公里 距西安北站约53公里。西安方向游客延西宝高速、行驶至兴平出口进入104省道向西延省道行驶约11公里到达马嵬驿景区。交警提示：前往马嵬驿游客行径兴平市区 避开市区道路。国庆期间每日下午14时兴平交警大队对马嵬驿景区进行交通管制 禁止所有车辆进入。　　8、咸阳乾陵 位于乾县城北6公里的梁山上 距离咸阳46公里、西安78公里 从西安可上福银高速、312国道前往 道路畅通 沿路有交通提示牌。　　9、咸阳袁家村 位于礼泉县城东北约17公里 距离咸阳26公里 距离西安50公里。从西安出发沿福银高速从兴平昭陵出口出 向北沿旅游路直达袁家村 路况良好。从礼泉出发沿关中环线向东直达袁家村 路况良好。　　10、咸阳汉阳陵 位于咸阳市渭城区正阳街道办事处辖区 距离咸阳国际机场10公里 从咸阳市区走兰池大道由40-50分钟车程即到。从西安上老机场高速专用线 过收费站向西2公里即到。　　交警提示：该路段为双向两车道 路面较窄 强过往司机低速、谨慎驾驶。　　11、咸阳博物馆 位于咸阳市渭城区中山街53号 距离西安20余公里。西安火车站：39路(南线)西咸快客直达；西安咸阳机场：机场大巴到咸阳北门口十字下车步行10分钟；西安汉城路到咸阳：59路；地铁1号线到后围寨：13路咸阳北门口十字下车步行10分钟。　　交警提示：咸阳博物馆位于中山街老城区 道路狭窄 停车泊位相对紧张 重大节假日早8时至10时 游客较多 建议错时出行。　　12、富平习仲勋陵园：位于渭南富平县城西北3.5公里处 距西安70公里。从西安出发 沿京昆高速到富平出口下高速 再沿荆山大道、怀德大街到习老陵园。若从富平县城出发 则沿桥山路至怀德大街到习老陵园。　　13、习仲勋故居：位于富平县淡村镇 距离县城5公里 距离西安70公里左右。从西安出发 沿京昆高速到富平出口下 再沿荆山大道到环城南路 到富淡路 习老故居。若从富平县城出发 则沿频阳路到环城南路、富淡路 到习老故居。　　特别提示：来者需带身份证；自驾车请不要超速 遇到暂时堵车 请不要插队 顺序通行。　　14、韩城市司马迁祠：该景区位于韩城市南部芝川镇东部。该景区距离最近的韩城市区13公里 距离西安200公里。路线：西安——西禹高速——芝川出口——马陵村——旅游路——司马迁祠景区；　　15、韩城党家村景区路线：党家村位于韩城市东北方向 距城区9公里 距西安约200多公里。　　路线：①西安——西禹高速——韩城高速出口向右——昝西公路——党家村。　　16、渭南华县少华山国家森林公园：少华山位于华县县城东南5公里处得秦岭北麓 距离西安约80公里。　　路线：(1)西安---华县(高速) 从连霍高速/G30 向东直行 到华县出口下 沿国道310方向 进入新秦路 沿新秦路行驶0.9公里 左转进入国道310 按照路标指示到达少华山国家森林公园。　　(2)西安---华县(低速) 从西安沿108国道往华县方向行驶 按照路牌指示到达少华山国家森林公园。特别提示：交警提醒各位驾驶员在山区道路行驶时 确保车况良好 注意减速慢性 注意对向车辆 注意避让行人。　　17、渭南华阴华山景区：华山景区离华阴市3.5公里；距离西安120公里。路线：从华阴市沿四十米大道至华岳路到华山景区；从西安出发沿连霍高速至华阴出口下 右拐(朝南)进去华岳路 到华山景区。　　交警提示：国庆期间 旅游景点迎来流量高峰 由于景区部分道路路面较窄 弯多坡陡 驾驶人应格外小心 注意减速慢行 不要强行超车、强行会车 尤其不要在弯道、陡坡停车。　　18、渭南合阳洽川景区：京昆高速西禹段：(距西安153公里)西安绕城高速——西禹高速——合阳出口下 经由洽川旅游专用公路(22公里)至洽川风景区。108国道：从西安出发途经临潼、渭南、大荔、澄县 经澄县寺前镇进入合阳辖区——合阳县城——合洽公路——福山——处女泉。景区公路驾车行经急弯坡陡 请减速慢行 注意观察 不要强行超车、强行会车。　　19、铜川照金革命根据地(香山景区)：G65包茂高速公路：由西安出发进入包茂高速公路向铜川方向行驶 约63.2公里后从铜川新区收费站驶出高速公路 后根据市内路线提示牌到达照金革命根据地(香山景区) 沿途可进入三原服务区进行休息。　　G65w延西高速公路：由西安出发进入延西高速公路向铜川方向行驶 约57.1公里后从铜川新区收费站驶出高速公路 后可根据市内路线提示牌或到铜川旅游服务中心咨询以到达照金革命根据地(香山景区) 沿途可进入三原服务区进行休息。　　20、铜川玉华宫景区：G65包茂高速公路：由西安出发进入包茂高速公路向铜川方向行驶 约101.6公里后从金锁关收费站驶出高速公路 后根据210国道路线提示牌到达玉华宫景区 沿途可进入三原服务区、铜川北进行休息。　　G65w延西高速公路：由西安出发进入延西高速公路向铜川方向行驶 约109公里后从玉华宫收费站驶出高速公路 后根据提示牌到达玉华宫景区 沿途可进入三原服务区、耀州服务区进行休息。　　21、铜川陈炉古镇景区：G65包茂高速公路：从西安沿包茂高速行驶约100公里到铜川川口立交下 右转过桥后向左直行约500向右 沿涵洞口宜上线前往即到。　　22、黄帝陵景区：黄帝陵景区位于延安市黄陵县 北距延安162公里 南距西安165公里 高速公路可直达。延安交警提醒您：高速公路行驶时驾驶座及乘客要系好安全带 不要频繁变道 切忌不可超速行驶。　　23、黄陵周边景区：距西安165公里 黄陵县国家森林公园、黄陵轩辕养生谷、黄陵万安禅院等旅游景点 景区道路狭窄、坡陡弯急。黄陵交警温馨提示：驾驶员要靠右行驶 留意沿线警告标识 行至转弯路段要提前减速慢行、鸣笛 遇对方来车主动避让 严禁强超抢会 防止刮蹭翻坠事故。　　24、延安壶口景区：距约西安330公里 从西安出发沿G65包茂高速??G22青兰高速??壶口出口下。　　25、汉中黎坪景区：位于汉中市南郑县。西安至黎坪景区350公里 高速公路280公里 景区道路70公里。路线：沿京昆高速西安?汉中中央大道?南郑?黎坪景区。前往黎坪景区道路为山区道路 路狭坡陡弯多弯急 且多临崖临水。交警提示：行车时要注意保持车距 控制车速。　　26、延安九吾山景区：志丹县九吾山景区道路狭窄、林木茂盛、视距不良 驾车要靠右行驶 降低车速 行至转弯路段要提前鸣笛 严禁驶入对向车道 防止发生碰撞事故。　　27、延安石门峡景区：前往石门峡漂流有两条路径 经304线(白马滩至大岭)、钟赵路(黄龙—柏峪—白马滩)即可到达。黄龙－柏峪路段。该景区道路改建即将完工 游客流量将剧增 可能导致道路拥堵和交通事故增多。目前该路段大车禁行 小车行使时注意保持好车距、车速 特别是超车、交会时 请先仔细确认前方路况 再行超车；会车时应减速缓行 避免因车速过快 转向过大占用对向车道而发生碰撞。白马滩至大岭路段多为临崖险滩 山体松垮 路面损毁严重 过往车辆需保持车距 减速慢行。　　28、安康岚皋县南宫山：位于安康市岚皋县东部 东起岚、平县界 西起柴垭子、岚河响水沟口 南临岚河 北至溢河。来往南宫山的西安自驾游客可通过西康高速抵达安康 全程195公里 然后沿S207安岚二级路行驶95公里抵达南宫山森林公园。从岚皋城区沿207省道至南宫山北大门到达景区约22公里 从岚皋县城沿207省道到南宫山南大门约24公里。　　29、安康岚皋县神河源景区：从岚皋县城沿岚城公路至神河源景区约51公里 从神河源景区到千层河景区再行驶13公里。另：从城区蔡垭沿月石公路、石横公路到达千层河景区约55公里。　　30、安康石泉中坝大峡谷：西安至石泉中坝大峡谷自驾游游客可通过西汉高速到石泉出口下 过大河坝收费站沿210过道 经过两河镇可到石泉县城 全程233公里。　　31、安康石泉子午银滩：西安至石泉子午银滩的自驾游游客可通过G5京昆高速南行150公里至石泉/佛坪出口下高速南行5公里可到达子午银滩。景区道路临江临崖 路窄弯急 容易堵塞 驾驶员需谨慎驾驶。　　31、平利县八仙镇天书峡景区：207省道(安镇路)——170公里+900米 距县城70公里 207省道传境而过 位于西安-安康-南宫山-千家坪-小三峡的旅游黄金线上。　　32、红碱涝景区：位于陕蒙交界处 距离榆林城区约90公里 距离西安约670公里 从西安驾车进入包茂高速 在红碱涝出口下高速即可。　　33、红石峡、镇北台景点：位于二里半向北3公里处 景点内设有停车位 可满足游客停车需求(节假日期间会增设临时停车位)。路线：红石峡、镇北台距榆林城区约5公里路程 距西安约576公里。由榆靖高速路口向东至迎宾大道与长城路十字左转 向北途径长城北路约3公里路程可达景点。城区游客可乘坐11路、3路公交车至镇北台站下车。　　五、自驾出行安全提示　　1、自驾出行请合理安排时间、规划出行线路 避免集中出行。出行前要通过网络、交警部门官方微博、微信平台详细了解出行线路交通流量预测及绕行分流路线 要提前掌握出行沿途服务区、加油站、卫生间分布及景区周边停车场分布情况 避免盲目出行 影响出游心情。　　2、自驾出行请保证充足睡眠 合理安排行程 注意劳逸结合 避免时间紧凑超速赶路 尽量安排轮流驾驶 避开午后和夜间行车 驾车途中要及时休息。连续驾驶不超过4小时 停车休息不少于20分钟。若感觉困倦、状态不佳 请选择安全地点停车休息 切莫在高速公路上随意停车。　　3、驾驶过程中全车司乘人员要全程系好安全带。驾车带儿童出行时 请为儿童选用适合其年龄、体重的儿童安全座椅 一定要避免怀抱儿童或让儿童坐在副驾驶位置。驾车时不要接打电话 不要边开车边设置导航等设备。临近目的地时要注意道路指示标志 路段不熟 或者不能准确判断出口时可以就近驶出收费站 询问收费站工作人员后再选择合理路线行驶。　　4、高速路上随意停车极易引发二次事故。车辆在高速公路上发生故障或交通事故 要立即开启危险报警闪光灯 在来车方向150米处摆放警告标志 车上人员迅速撤离至护栏外安全地点 打电话报警等待救援。　　5、驾车行经农村、山区公路要谨慎驾驶 夜间驾车要减速慢行 注意观察道路情况和交叉口车辆、行人出入情况 与前车保持安全车距 切莫超速、逆行、违法占道行驶。　　6、上高速前细查装备。俗话说“在家千日好 出门一日难” 开车上路 特别是上高速路 一定要提前检查车辆和“装备” 以备不时之需。机动车上高速公路行驶前 最基本的检查有七项 包括：轮胎、燃料、润滑油、制动器、灯光、灭火器具、反光的故障车警告标志 并要保证齐全有效。　　7、保持安全车速行驶 切忌车速过高。在高速路行车最重要的是保持安全车速 不可超过限速标志牌所限制的车速。　　8、高速行车最忌讳的就是动作生硬 转向时方向盘打得过快 角度过大都可能使后轮失去抓地力而导致车辆失控。当前方出现意外时 不能手忙脚乱地猛打方向 应该在减速的同时尽量舒畅地转动方向 让车平顺地躲避险情。　　9、掌握制动减速的窍门。先轻踏制动踏板告知后车 然后再减速；要采用间断式的“点刹” 以防车轮抱死打滑(有ABS系统的车例外)。　　10、驾驶员朋友们 您在出行前请提前规划好出行路线 注意高速公路出口提示牌 以免错过高速公路出口 如果错过可从下一个高速公路出口驶出 切勿在高速公路上倒车、掉头、逆行。|http://www.shx.chinanews.com/news/2015/1001/42260.html|2015-10-01
其他媒体|2040013687|zhidao_baidu|电脑/网络 > 笔记本电脑|ZHO|2015-10-01 15:11:01|东风悦达起亚k3多24期0利息是真的吗|汽车|http://zhidao.baidu.com/question/626524537027364924.html?fr=qlquick&entry=qb_list_default|2015-10-01
各大媒体|2040368697|qc188|车主说车 > 紧凑型车|ZHO|2015-10-01 18:32:02|绝对的高颜值 朗动6000公里用车感受谈|本人生在一个小地方 普通的上班族 本来没有买车的想法 去年3月份和朋友一起考了驾照 5月份就拿到手了 看到身边的同事一个个都买了车 再加上几年工作有了点积蓄 于是乎就产生了买车的念头 每天像吸毒一样 关注这每一款车 无论几万到几百万的 几乎天天看 其实我对车蛮了解的 因为我就在本地的龙头企业“东风悦达起亚汽车有限公司”上班 所以比一般人接触的多 本来想买公司里的K3 公司还有员工优惠 但在盐城k3的太多了 再加上每天都要面对它 有点审美疲劳 正好今年车市不好 其他品牌优惠都比较大 于是就开始关注其他品牌的产品 价格和k3差不多就好了 当时心中有几个目标。 ————————————————————————比克的新英朗是第一个看上的 漂亮和内饰都不错 但因为当时优惠少 就放弃了。 ————————————————————————大众的宝来是朋友介绍的 本来对神车无爱 但老爹喜欢 说牌子响 不会太掉价 去4s店看看还是无法接受套娃的样子 果断放弃。 ————————————————————————吉利的博瑞 一款非常好的B级国产车 高颜值的外表 超高的配置 空间也大 当时很想买 但因为才上市 本地4s店连展车都没有 下单订车 不知道要到猴年马月 只能放弃  ————————————————————————北京现代的朗动 其实这车一上市就很喜欢 但当时驾照都没有 再次关注起 还是朋友介绍的 自己居然把它给忘了 知道朗动和k3是亲兄弟 所以我也没有太多了解它 就去了4s店 要求试驾 然后就是和销售顾问一阵唇枪舌战 最终优惠2万 送脚垫 车膜 和一堆不值钱的东西 在这里说一下 我定的是自动领先版 外加选装包 落地12多。 好了不多说了 开始上图 照片都是肾6拍的 拍的不好大家见谅。 ---------------------------------------------------------------------------------------------------------------------------------------------------- 正面来一张 牌照就不挡不 有盐城的朋友看到打个招呼。 45度角 就是车头短了。 开门的侧面。 很喜欢这张 led日间行车灯 没k3的霸气 很喜欢侧面  翼子板 还蛮硬的 再来一张由前往后的 右边  车门 厚重感不足呀 门把手 带无钥匙进入 喝茅台的嘴 17寸大脚 北京现代 伊兰特 带折叠的后视镜 贴的防全景天窗膜 后屁股 网上买的后唇 大灯特写 尾灯特写 外面装的迎宾灯 感觉不怎么好看 后装的无骨雨刷 一片狼藉的后备箱 中控全景 用料不错 很多软塑料 放杯子的地方 无视口香糖 扶手箱   [1] [2] [下一页]|http://www.qc188.com/czsc/201510/127066.html|2015-10-01
其他媒体|2040474586|zhidao_baidu|生活 > 购物|ZHO|2015-10-01 19:34:01|起亚k3飞歌dvd导航仪倒车影视没用是什么问题|硬件|http://zhidao.baidu.com/question/938769346180125452.html?fr=qlquick&entry=qb_list_default|2015-10-01
기타|2081878669|xincheping|首页 > 讨论区 > 购车问题|ZHO|2015-10-25 18:07:12|落地10万 自主车和合资车相比 谁更有竞争力？|由于手上预算有限 只能买落地十万以内的车 想请问一下自主一线的品牌像艾瑞泽7 逸动 帝豪 悦翔v7等车型 这些车型的产品力是否跟日韩系的的像朗动 k3 卡罗拉 雷凌等的车型已经差不多了呢？|http://daogou.xincheping.com/115007.html|2015-10-25
其他媒体|2082017101|difang CN|地方频道 > 滚动读报|ZHO|2015-10-25 20:00:01|期待在家门口赛出最佳成绩|2015ctcc中国房车锦标赛（盐城站）将于今天11:30举行发车仪式 标志着中国最顶级房车赛事的超级量产车组、超级杯组、中国量产车组等3个组别的比赛正式开始。史翠英群星车队剑指盐城橙色军团史翠英群星车队在上海佘山第三站取得5分后一直蓄势待发 这次终于重返ctcc赛场 盐城晚报记者昨天在赛场内看到 史翠英群星车队的招牌非常醒目。由于战略调整等原因 史翠英群星车队在今年的参赛场数较少 但这并没有影响车队的整体水平 这次 该车队以俱乐部车队的身份参加ctcc超级量产车组。去年 史翠英群星车队就在盐城有着不错的发挥 两辆赛车都取得了积分 并夺得了俱乐部杯年度总冠军。科鲁兹掀背的赛车经过多次升级后取得了很好的口碑 而赛车的实际表现也证明 车队的付出是值得的。老将陆淦表示：“每一场比赛机会都很难得 无论是我还是车队都会珍惜这次比赛。在试车中我发现赛车的整体感觉比去年在盐城站的时候好多了。我们将全力以赴 为下一个俱乐部杯冠军而努力。”北京现代担忧车重影响发挥北京现代纵横车队再次登陆盐城街道赛 去年 北京现代曾在盐城年度封王 夺得中国量产车组别年度厂商杯的总冠军 车手崔岳也摘下年度车手总冠军。可以说 盐城对于该车队来说确实是一个福地。目前 在中国量产车组中 北京现代纵横车队暂列第二位 现在遇到的最大挑战是规则加重上 因为崔岳处于车手积分榜的领先位置 而他的赛车又是全场最重。在盐城这样需要出弯加速度的赛道 赛车上每多一分重量都会降低速度。虽然车重令崔岳比赛形势不利 但他表示会与队友一同在盐城街道赛上做出战术配合 争取获得更好的成绩 “我们的赛车速度还不错 但是比去年慢了一些 目前试车结果还可以 车队还在努力寻找适合的调校 我和车队技术人员一定会克服这个问题。”东风悦达起亚与k3s齐发力ctcc上一站在上海国际赛车场进行 在超级量产车组中 东风悦达起亚车队的叶弘历斩获生涯首个ctcc冠军奖杯 东风本田车队的谢欣哲与何伟权包揽二三位。叶弘历今年是首度加盟ctcc厂商车队 参加全年的比赛 此役 叶弘历终于圆了在ctcc站上最高领奖台的梦。比赛总共10圈 他凭借完美的发车超到了第一位 之后虽然跟何伟权互有过招 最终还是顺利第一位冲线。叶弘历证明的不仅是自己 也证明了东风悦达起亚与k3s赛车的实力。据了解 这台k3s搭载的是韩国本部研究所研发的1.6t发动机 以量产伽玛发动机为基础 瞬间可以爆发出300匹马力 缸内直喷和双可变气门正时技术并重 扭矩更高 耗油更少。为了应对不同赛道的艰难考验 东风悦达起亚技术团队还对底盘和悬挂系统做了针对性的校对 为车手打造了一台极具操控的速度战车。盐城晚报记者曹恒锋|http://difang.gmw.cn/newspaper/2015-10/25/content_109648732.htm|2015-10-25
기타|2093136331|ngzb|新闻互动|ZHO|2015-10-31 23:11:01|广西女诗人陆艳辉获“中国青年诗人奖” 获奖作品：《心中的灰熊》|"马上注册 结交更多好友 享用更多功能 让你轻松玩转南宁您需要 登录 才可以下载或查看 没有帐号？立即注册  x       南国早报网讯    据新湖南客户端消息 10月30日 首届中国青年诗会在湖南湘西自治州举行 诗人黄明祥、陆艳辉（女 广西）、晴朗李寒获得“青年文学•中国青年诗人奖”。"" S: @: r1 v# ]6 h; }8 ^' k4 F7 l6  ! m( Z. P中国青年诗会由著名文学期刊《青年文学》发起和主办 今年是首届 今后拟每年举办一届。该项活动以“发现、培养和推举新人”为宗旨和艺己任 每年遴选在《青年文学》“汉诗”栏目发表作品的优秀青年诗人参加 通过“作品评奖和研讨、社会实践和调查 实地采风和走访等丰富多采的形式 展现青年诗人的创作实力。”- {  Q8 s  S9 B5 [/ M9 M3 _0 h/ T; r"" r8 m7 x% y中国作家协会副主席、书记处书记吉狄马加从北京发来贺信。他在贺信中表示 中国新诗将历经百年 对新诗的回顾、梳理、展望 和对脱颖而出的诗坛信任的提携表彰 都是中国新诗蓬勃发展的原动力。鼓励诗人创造出更优秀的作品。"" o/ w8 l6 e% A5 ^0 U: x| _5 Y. J3 u9 K0 K诗人陆辉艳的作品《心中的灰熊》、诗人晴朗李寒的作品《月光下的磨刀人》、诗人黄明祥的作品《从未有人走过》获奖。0 w& y0 u0 j6 e- OQQ图片*************9.png (868.15 KB| 下载次数: 2)下载附件 保存到相册16 分钟前 上传4 @3 B( i  B+ \. Y& s 诗人陆辉艳。7 y"" A3 y| F# c4 A  G5 L3 Y$ P- Q0 D. c获奖作品 ! j: a) m+ `2 F8 [2 x( F/ G- ~; D7 f8 s一、陆辉艳《心中的灰熊》 7 O0 [1 `* s: Q2 b' Y+ R"" V2 ^# n& w; X/ S3 ^8 _| G/ N- p; C# Q6 S1、反 面- u# @- I9 P/ Q6 C8 Y"" D3 C& q- Q$ H+ \5 D3 B' o/ \9 L& N6 G"" C& ^7 e* ]' E那是个诗人。他们说 但她不喜欢交谈! s' \- g3 F7 L8 v9 e1 j- G3 ]| A' E* c8 u! ]! _"" V3 G4 [3 N- h5  : \' [7 p& i! z| q9 l她避开各种形状的镜子 水泊 大理石 一切) o% @' j6 u* [: i  l( Y3 g; O"" A4 g0 H2 u0 m(  . h2 Q) ]# }8 q; W  X4 k& R反光的地方。它们映照或遮蔽大地的秘密1 A# s- G2 `) y/ Q# q/ r4 h: R4 ~) q( F! o  y' p# R) T9 p- v7  ) U0 o+ \相对于判断 显得力不从心| z! ?  I8 Q- g"" l0 t: Q5 P+ G1 d7 b) e! c) I$ d9 q3 s8 Q$ ~8 ?# K7 g7 X9 H她穿平跟鞋赶路 像一阵稍纵即逝的风7 Q7 Z! z5 z| `:  &  4 Q/ P2 Z9 k: [) N: V/ o| p/ @  i8 T1 ^9 o1 i9 r' q但在穿衣镜的反面 她遇见了# @| x) R+ ~# k: H4 R: Q| ~( I7 R5 I+ }. o* F* o| h荒草般的自己 她甩一甩脑袋% K3 a# b) s8 }* g- V; D9 f4 O$ y/ N% ^4 P& c: A1 ~' N( s. d8 l8 Z& C9 p' I' F# o第二天去了理发厅3 _# _7  6 U' v5 _5 i  S9 D2 M' A  \! W9 B: u/ ~' F/ H/ H在那面光洁的圆镜前"" K- E1 T! q* w$ o& h2 r9 k/ h5 S- j| H9 X. X4 j) d% J她紧闭双眼 让造型师把头发$ J/ F0 q. {9 U; J  G' g7 }' C* r3 C; z3 I0 I"" D# [/ z& x$ T9 `0 e- l8 j弄成了蛋卷状。隐约 她听见9 ^  t! m- ~* v3 x1 {& g0 n. v& h# s! h# t! _| D"" ^6 B/ I. `% w! H| Z; _6 v蛋壳碎裂的声音% X& J+ G3 G9 l  Q| I- U2 y$ @8 s! t* k4 g( r! r% e$ u8 M| p她踩着脑中的那些碎片 上了204路公交车; d7 d8 l% y4 K  D/ s/ _4 d5 z5 o4 Z& Z. f) g5 H2 b7 ~# p- S2 F* b% r; F一只手抓住铁环 在发酵的人群中- f/ t$ Z/ _- T6 t0 C7 A7 L2 ["" c1 F  I3 ]+ H% H0 i/ `2 H"" m6 o5 @: M昏昏欲睡 错过了站! b7 w+ `7 p# H% b& p+ i7 `/ x* M5 z0 p( n( J9 Y8 @' K! L' Z( V"" _! F5 R$ h( H9 x当她抬头 黑色窗玻璃上映出法令纹' o$ X! I* T! ^! U* A6 `% E3 y' Y+ k* t$ D. n& k3 I2 c2 v&  2 _6 l多么深的时间的沟壑 紧攫住她的额头$ t: v: R1 }; S2 e$ b( c( ^% A' u4 J  h5 t+ T2 B. K/ p6  3 k! i3 a对此她并不介意。扭过头 下车5 V. b/ A+ N7 p1 c: q6 J# \) n0 ]# A) {; @! E4 ^1 z* I' ^( V( S8 X泵入下午的热浪――带着她的新发型"" Z+ e- i& u- A. E4 @4 S& G7 f) c+ @: i: k- D& n3 d$ X3 w6 l3 ^2、只差一步' \: J: L- }0 w1 Y7 n"" [6 k% R% _- d- e. k9  - F| ]# T#  * {; r2 L那是一道闪电的开始。阳光的移动  f"" f8 [0 M$ t4 _; h* ^"" O2 h5 l; h; O! T. N6 A  D. A# b7 ]9 Z制造了一片槐树阴影。跳探戈的女人: x&  4 l6 ~6  . ^6 ?!  ; n# N2 e1 V) ^6 z! C& j0 C6 M双脚钉在大地上$ R! P$ E0 ^3 k/ l8 C1 R* N& ~6 j3 x# K; o+ A"" n' p& Y9 u( i( V#  她表情严肃 仿佛另一个人贴紧她的脸; s/ ~! ^/ q8 P) {3 }& [% T9 W# o+ ?0 ~; ?% Q' ~) s$ L| F0 C! K8 ^3 y+ ^/ E4 ~& Z6 j; Y追逐、躲藏、踢腿、腾跃、270度旋转4 A. v8 `6 C8 ~& c! `+ ]0 v& u( {- b0 X; m"" s9 T% ?  v# H. o  t9 s. r8 I0 i0 \# j$ \7 y""  9 m/ T――她搂着一个不存在的舞伴! ?+ Q% ^/ {' c5 Y3 D4 W& R6 _' E  x/ u) c| ~'  ) R# V1 \9 x)  ' b; b在一个断音处 她突然停顿。像是一幅剪影|  $ O- u5 h1 I$ @  F9 K: l"" e% z2 m% H*  7 R| O; g( k! u7 k8 p一幅未完成的雕塑。望着空荡的前方& b* W) X! {2 j2 `5 `- g/ ?9 p3 Y5 s' a  ~5 g1 f! i: t; n! c% O3 G/ O9 e) c似乎在等待下一段旋律  M$ H"" C. o- M* e) R7 k; L6 l6 o6 H7 v( y0 _/ d+ W8 l% d8 S$ S2 h- C+ R1 ^' B! D或者未出现的人/ A' a: z8 M+ f4 J; j) W% R$ z( l6 ]9 \* {$ ]2 l) }2 I- V; V  K) E7 N& y后来她深吸一口气 开始东张西望% p0 r"" D) \6 g   4 o8 L! W# q6 F% m1 d3 s& I+ h; y"" ?9 [: b8 j1 q| m: F* p8 @像是提防秘密被人发现1 H/ H1 d/ x$ N( F/ }! N* ^& P* L. ^8 f+ I+ r! q5 x1 a. P  e6 L; `7 s| A6 G5 s# b我听见黄昏咔嗒一声+ D  A| e5 P+ w2 M: O% ^0 Z: `; T% J$ [  T1 T5 k( h/ p5 k8 c  T9 j* M舞曲仍在循环播放：只差一步。' G"" o6 t+ B/ P| z| ^7 n' L. e7 s7 U; l( _. B- ]9 P; Z1 W- S只差一步。尚嫌不够。永远是这样- Q"" k' s2 P9 A- h- B! Q( ]9 c2 T1 D5  % B6 O5 {2 N| p( d) S2 X. d2 A3、力 量% w- Y! Y' G3 r8 o/ }9 _  [* d/ w( W5 a% {/ E! h( B"" J7 m' A3 ~$ X  C. S% A- X那看似微弱的 胜过一切5 `5 W/ b| Y3 H| s. P) p3 y! z3 D  L# j6 C| Q: g) N1 ]4 X' Z) I$ d种子顶开玻璃瓶塞9 n( N* y* Q% A6 s3 F6 ^& \5 V9 e$ h7 q% K1 L1 Z/ c& X$ r蚂蚁抬着一块面包过了桥| D4 q. G0 Z9 [8 o( G0 b7 ^- i( E4 B' m4 I/ D; N# l+ }| A  J+ T4 a: E4 p- a羔羊眼里流出泪水( g| r0 N2 K9 v3 ^$ l:  8 q0 ^% s8 u5 _6 L0 }9 w4 ^# ?4 N3 `| z# {* X它将人类弑母羊的刀子藏于自己身下' C6 {3 @0 y* i) _( X2 c& R2 H- O9 \| A' W! t* Y9 i( j- e+ m( g/ s( L: ^: G; s$ I黑色枪口对准一个手无寸铁的男孩9 [. g7 ^6 A2 o4 _6 {; d1 H8 b| L7 _+ i% R) n  k: A) y"" y. X: N1 `; h0 k他把鲜花插在枪口上| l. G"" E# s; x% M!  ! X| M"" a( D7 u( ]+ Y+ @4 ~$ P'  8 O: h4、然 而/ w| u. L& G9 D+ K* P7 l1 G5 P& \| a' O! u8 _$ w9 t# w9 n& B  X6 d0 K0 c7 ~陷在凌晨的腋下;马匹站着酣睡。5 Y6 ?! H| r( ["" M; S4 G+ Y| O+ z( Q: X2 }1 ~% \1 j' ^7 `# f1 s  w那洗盘子的女人 有湿漉漉的手和孤独。# j1 Z0 w5 G( K1 G| `| o* R5 j| H) \; v3 X9 @' n9 g  y0 w0 K0 x/ d0 U0 w她听见盘子碎裂 时间的胎位移动。"" ]"" R7 g5 q'  5 G: n9 U( r3 r' h; U! q6 S( Z& ^+ Y4 V0 s; d4 x. L( S我们头朝下 星空广阔 在下2 I* H+ v; ]4 s& ?' ?# b"" Z8 C4 L3 t2 m/ t  O) F! x1 d  i  x; T抑制不住猜想这些时 她的脸部绯红- N4 }. u2 r; p( L% \& q; t| W1 r( j4 h"" F6 Y3 }6 }5 {; H; K) a她想用故乡的语言去纠正那些本地马% Z"" _' z! S3 i% E1 z5 m- @2 N3 F- x( ~! {+ t  U5 N3 ?2 @) X4 ]5 X可倒春寒使喉腔冷却。1 b* @6 S  m"" ?6 f2 F! e$ g3 n! Y8 f. W) U/ G( Z% d% p+ `8 U5 \& ~9 Y. \( b昆虫们集体在清明前噤声8 k5 k4 r7 i0 S1 d1 H5 s( Y% ^; J* q| n* f% L3 `) _( M! d- H: I5 s+ W* c! g1 k! i# Y: Y' \* p& X$ x5 O所有的夜晚都集中到这儿  O* j"" n/ q7 o"" _& G"" G9 h: b- M- `/ d' Q9 G| }+ a( n$ X; o5 C# m"" E# j/ I* ]2 _然而她还嫌不够。桃树已经结出桃子9 R2 b# K# t6 ~; x& F3 w2 q5 M( I5 O+ G$ O  r8 ^* o- o9 e| v* b- B- }等到五月 人类把它们摘走 鸟雀会不够吃5 {& P6 I# A+ l9 j# @& `8 I4 @5  3 O. [9 W8 F* D- M9 v( Y不是没有可能 打开山中屋宇$ g2 ]9 Z3 a) e! u  S"" s( z+ @: u3 U! v| F| R# ]2 n) U- f. I. Q- _8 I. S6 ^+ Q) o天边的鱼肚白会蹿进来 长住6 F# ?. _! D* D$ f$ _9 A0 D3 H+ B2 d2 C4 P8 e( b  T6 U/ n6 _( f) b0 N/ q& U( ?1 _蝙蝠像黑色的文件夹 倒挂着合拢& ?6 b* d3 Q& R) l2 H/ E5 K# f* I1 j$ p8 h- c; _! M( b0 E4 i! j- B! w' @* T然而只过了一刻 她便倒头睡去4 V0 W- n) c6 d$ Z3 G5 X- D"" o% B3 F/ A5 B! G) T.  $ ^' j9 P+ h- A: \+ S在未洗完盘子的长凳旁$ s+ J/ G% h) B+ \# r7 X# @8 g. L( X4 @3 T' {. p. w! T1 j- y4 J5、搬 离' y8 Y| s& x. o/ M% [3 B0 j/ k: z7 C8 J# X- s& o% H7 {"" }* M& ]0 K( }他们搬走了你的桌子、口盅和文件4 p5 b( I$ A8 G7 _  s3 Q3 S* U2 L6 _% i) J8 J) y(  $ V) L"" g4 E1 o: C$ o2 H"" S3 J水养的绿萝也被倒掉水4 e9 z3 Q. F* j/ c' a& J( U$ I0 q! d2 {0 `|  $ L$ B) s装进一个塑料袋里 连同背电脑的8 A"" v+ I) L| f0 R- r# c  r5 d8 Y& l$ O- ~7 A- N0 v| w8 b+ o! x工人一起离开。你看着腾空的办公室5 p* Z2 S* h) G; p( Z% F4 Y% v0 k8 g$ n* g) [! l4 b  e7 ^; n2 X; _4 I不知该说点儿什么。下午的阳光) _; O% V/ x&  2 l- M* v- g. ?; g. _3 u& N3 P9 q& p% g) ?! }从后窗爬进来。满是灰尘的地面/ j"" m| k- j5  . M$ }. `| x1 L3 G3 z+ H' `4 i  D& a: S4 r! b# F| ^# [( Q被照亮。你竟然与这些尘土7 d5 e1 R( J2 t1 g! _3 w; e  O+ c# K9 @) ~8 e3 S& L8 F4 A7 U* l% v. D| G4 Z2 m- w! q相安无事地共存多年而无察觉  x! u+ n' e8 L) T* g9 J4 @! [| P! U"" J7 `- R; F"" R+ a7 b0 X  ^5 `8 K它们被太多东西遮蔽 直到有一天! U- o! N7 f9 _5 F) q/ j/ v  I$ p7 K"" z# P+ e+ E* e! F' e- R6 z9 `- t! S7 C- A& C无辜地显露在阳光下。你将抛弃它们: i: M/ r$ l8 h1 ~0 \( [4  8 J0 E2 M. [* h9 a1 \| }  T5 Z3 [3 H1 u5 f. L5 z到新的地方 继续耗费你的光阴 激情( C: n$ z+ ?/ I$ e& O2 _7 i; [& j* l; t9 T* M& D5 E3 P血质的孤独。你需要这样。你的同事0 g* H! O; _+ Z& @- f6 V* V/ }# U| `7 c# F) V: Y7 p/ z) W| \0 ~% m. [8 b9 a在对面新装修的大楼走廊上2 Q; ?: }( n( Y| s3 p& q3 G2 B3 b2 q- s7 s/ B: {- }6 D/ M7 \' K|  5 G. }"" h1 f0 k+ I9 K笑着向你招手。你关上窗 但没能9 V. T"" b"" k0 O& y) r) w8 e8 K2 g7 z"" v! r0 v  ?6 }5 V| e% f2 j0 R5 z| R. q关住阳光。帘子已被拆走7 g& x( m) k# O: C' ^5 S3 f. G"" [. m6 S- x  q7 t& t1 E0 Q. w- g3 x5 o1 {像每一次的搬迁 你抱着你的物件"" m6 L$ Q0 d& A* m. L: P4 \% E6 i' z| v. X9 A4 x& i0 [6 N% C. U4 m. s' T' Y6 M最后看一眼那个有你气息的地方& j5 H4 {9 A  d' ^- r! k- T9 a! l1  4 W6 z0 X8 z- J#  ; {# e( \走出去 反锁好这道门| `; y8 A  ?8 v4 V| ~; ]1 A6 v* {! C. D5 c6 I3 S' ^8 ?& O/ H7 u5 c& y把钥匙交给另外的人# J- v& G3 a: ^0 W7 u* b6 O- A( x3 J. q! V# Z3 Z"" Y5 m6、叙 述8 E"" G. k. ~5 Z! o2 g- V"" X( S- Q5 z2 S9 e! ^/ K3 D-  ! Q; H* gY 我乐意向你叙述 一天傍晚' w- P7 }' h# e% {| l8 ~+ T7 l' n' E+ m6 Y+ v+ R3 r/ X4 y7 s6 v"" Q- p) Q- e2 [我是怎样走在江边 看茫茫夕阳"" t) Q: L# B; @7 ^9 f$ A0 A# I& U+ n*  | }0  2 z0 b! P' t6 D落下寂寥人间 江两岸的人们! r! ^: E: O% Y1 R& u0 o   9 r! L; a/ A) G0 f  y) G$ T5 w纷纷收拾工具 离开田间 回到4 l' O9 E8 N6 f0 V! f' t  q0  ' V"" I9 s- @# _1 l: q/ j0 i9 r% S' e# M2 E9 A家中 生火 做饭 升起炊烟  C5 T- x# q3 w1 W; ~  z| y  B. _5 \. }7 u: G! p) B(  9 H; e| {/ l+ g我曾低下头来 看脚下的石子! b* i8 C2 n$ d$ m- L- u2 z7 n% I- O& U- P* z; A1 D% l0 }7 b4 o"" g; O多少年的洪水 没有冲走它们* u0 i7 H(  ) v1  * _) Q# E)  . l6 r| U1 r0 t3 o+ Z0 g2 x  [# y2 R7 [1 Z5 W+ k: K) I: H3 w& U光滑 圆润 它们依然在这里 陪我说话* Q( [4 a) Y2 j2 z- s* y) h% R$ ]: K$ K2 K1 I| H| Y: D: b. {看天上闲云。因为喜悦 而将手停于1 j$ x3 r& {( N"" d  M; n: M. f5 L1 U& \0 m; H: Z: X3 y0 E1 C' D/ [0 o腹部 听到里面传来原始的搏动& o4 V: z+ e! p. z"" j/ h| G. `% v  W9 p) ]1 b; ~( g3 [的确 我不知道的事情 正一件件发生$ v+ O7 W5 y| a0 _1 E4 v. u- z: t6 d4 m4 ?% }/ O2 ?- Y( x0 ^  N. K! ]% x比如一个小东西 正在我体内生长- W8 i) w% N0 L! K# ~6 X7 j2 b1 C4 a9 {+ @( A0 }+ o* \| ~- D2 i5 H. o' z像个胚芽 圆形 走动时有空旷的回音6 O| M$ ?  A6 \2 [2 a0 s* w: p) g) o% ]| A+ [* q' o+ Q% w8 D' S5 i+ H# X4 j) \   ) Y$ h  m我承认自己固执己见 必须为决定) ^' {0 I| l. J$ U1 g2 T7 R  K& h) k5 ^3 b! e3 b7 j/ q$ q6 f& L"" z/ z$ l7 J承受一切：放下人世间的享乐* U7 x& h+ B# T: C7 I. C+ y% W% ^- y& P9 \| U9 t( }. D6 T1 y2 A% L% m像闲云般散淡。必须俯下身来1 w6 c; v8 Y' J9 V4 M0 r/ j# T& q+ c! g& s: s5  "" Z! O( d  u. ^. q) X' H倾听大地的胎心 安静 秘而不宣) ~"" A$ h: d% X' W"" q# s* y0 J4 @: h: @7 }# z. k2 b+ P"" I/ n2 H4 M% H! f! X. a0 }有时我站在矮松林下 听到风吹拂: m' ~; \| @9 p- X; u0 [1 W- U* M8 A8 e6 q7 `| c松针的沙沙声。我知道了：这一生简单的智慧( Q- P0 ^"" N8 o| e0 H  J' i5 R3 U; e$ e3 C+ k; A9 d0 K* h3 n- ^. g8 A' b和简单的善 风一样的 用我的小半生1 X9 R2 q8 a1 C+ Z- o0 n; ?) s6 I$ E1 `- h3 P3 T| o# Q8 e+ w去明白 而用大半生去学习2 q| u; W2 P; U8 W5 I( {* J: V+ C| \5 m3 D0 B& v6 U! y| }+ p2 k' h0 A) o我自信还有足够的时间 因为上天给我的+ m; {4 V* u| ^( Y. F) ?* ~% L+ X) T7 s7 F9 r: K0 E8 j3 z#  0 R  Q& Z' _5 B  C+ ]4 y又一次光芒 它已经开始| T3 B- @9 m3 X| [: b7 p9 g( J; `/ }) c7 J| p! M+ Z8 X# V! Y3 b* J6 ]7、落 日"" L5 L/ J! P# `| J"" G% V$ Z5 S. c4 y# k: t! D: `+ T  k0 S$ X8 x% n落日绕远山 许多事物的影子) v8 l' ^4 Q"" N7 A9 _& v2 g+ O9 ~: }+ n- S; @  L- h& P! ^5 g8 ~在大地上浮现出来。在一块岩石上' X- d& c5 h! R7 G% t  v( e/ l: Q6 F% }3 v0 q/ Y% }. ]  M0 w| s0 t9 U"" p& e我们的手印和脚印 多么像是* `9 }0 T4 W/ g* \0 S' V| o1 c"" _6 x: p( ^5 I4 r0 I$ k0 Y9 @| m刻上去的。我藏在树的% h6 y0 b  r| }& O! U. F9 h% }% q; [5 Y! z2 S+ p/ k' Y"" Y& W6 I5 _阴影里 你看到我 仿佛我们 也像是8 b3 J0 ^6 a$ O9 ]0 S7 n4 o+ O1 v$ ~) v4 ~7 n- J) s$ O3 J. O3 ~7 @$ A# f# e: z刻在了岩石里 不会交谈3 U  O% m8 u' P5 r"" P:  7 I: I6 u1 N3 J2 F. `5 L"" I% H9 I* T% V2 ]' j也不会亲吻。但是当我们走得远一点儿) v: J7 M* W5 V* }; v) q) [& J  K& Q$ ~7 x* }( h"" o' v/ g7 O8 o落日就落在了我们身上: J% b7 h"" G; \/ A1 j7 ]7 r' L1 e. r"" t1 T9 w' _1 S8 Y& W' m- f/ ~* f时空弯曲 你几乎要质疑自己所见' p; E# h. }+ N1 r) F2 i' J' [! x2 k! M! ^/ x  Z6 K| D1 O6 L$ P/ }. I( o+ x! n像一个真理 像是一束光( E$ \: A9 I0 q: _; ^) ~  J  b# j- n0 Y( b. u  V* U4 p长期睡眠在岩石内部2 l0 f5 b"" N% f! {) o0 X| j* f$ v( M9 ?) Y- q| }9 M2 S6 C1 v8 O/ {6 i* n- K直到时间来拍它的脊背8 X# X| b| E- k5 T"" {8 g5 g& ?3 C  s! D- f"" J+ z% z+ v/ k3 M1 a  }) u8、心中的灰熊- f3 F% I7 B) y2 ~. F% O- w1 s9 D8 N3 M% a9 }8 @0 ]$ u. a9 _: w0 a"" @/ I浅睡在他心中的那只灰熊+ _1 D2 p& q8 y/ K! H"" y) L| M* k4 U3 S  t% q: `6 e3 W9  9 A. ]再次咆哮起来 扑向他。“在黑暗、隐蔽的9 w9 @3 R& q7 T% H& M0 K: p: `. ?# `6 W6 p& Q2 r* O! w8 v) C# L$ [. u地方。”这个声音使他发狂"" B2 F8 A) S. M; m/ \# w! e; E/ y2 n$ v| a/ k  ]8 M+ R) c# ?' r+ T& D6 D使他不顾一切冲向荒野$ C. f- M' }) o+ X| j6 r4 ?8 ]. `( ]0 C- {: w# a  t# i6 `8 j' @% C你握紧鼠标的手 也跟着他: q1 Z$ h8 R8 j% f7 x! V- A(  7 a0 n1 K4 Q% T+ z! j8 n"" {6 T3 M6 S! _在风中狂奔 因为激动汗水濡湿手心( z+ ]. K& e  X| }8 b5 y# s: B8 o+ k( E8 {! r6 J| D' ]"" [1 {  ~  c你按住暂停键 想让他: r# v0 T2 i) K* J# v/ c8 I"" J& S# y- i4 U& J"" a6 {8 t& }9 C2 Q& B不安歇的灵魂停一停 停在时间的某一刻4 i9 y! B; m; X' d. R6 i7 j% o- u. }' z$ Y| a! G6 V8 q(  * B7 O8 i"" J"" _% Z3 i9 }6 w- L但无异于企图熄灭一场蔓延的| {2 f' e% Z( ^7  ) @$ Q$ w0 ?4 S  x8 L3 n. Q4 P0 {8 u| u; p| w"" H9 s平原大火。你眼睁睁看着他% `"" l4 O; Q2 K$ C"" }: r8  | Q0 k"" N4 ^; E1 k+ l8 Q$ r$ l$ c+ K- z"" W在一部传奇中烧伤自己。他去牧马 去狩猎) u6 ~&  ; \: {0 }5 O| H8 p+ F' C9 J' j6 T5 R! P$ M| b! ^9 k) g+ n3 v% o% B生来听觉敏锐 能清楚地听见- V$ Q3 b3 C8 ]7 [' ?( q* _5 r/ j% I1 N* m  v| o# T  h"" q| e0  从内心的密林传来灰熊的声音* h. j: I+ ^"" {  g+ K. D# R( v5 H: M8 Z* D! o8 h3 C- l* S# H! @) T2 g: x; N自由的生命 如此放荡不羁- B/ B! S: c& ?+ i"" V- O| P4 j/ a+ U4 U) N3 G3 s' g. l. v5 y- M6 K"" }现在你将别人的经历一再扩大& }| [+ v( ]: W5 d9 ^6 O! h: q2 p6 l"" J| O' m* k. P- ]; _+ j3 M1 W)  8 E假装是你自己的一生. P: A2 i7 C/ K1 q% z% ~  d0 l; [4 I3 ?/ w+ ?7 `  X+ n)  "" G| ^0 H2 O# l% `2 b; U   以此安慰你那颗青春将尽( T  C. y5 B$ J2 a: v: i  j# j# `5 d5 a5 M4 I; x: n2 Z' o9 _: F2 {而不够勇敢的心 “将众人的明月 6 u( v9 v1 ]4 Q+ c  J/ W6 J5 i+ X) C. s* k+ e7 i/ C"" v! H/ m9 z占为己有……”& E) }$ g8 N| u+ A% _3 m0 i: `# ]6 Y7 `/ C# x* Z| Q& g: d+ N: A1 u4 e$ r为此你感到了羞愧 脸红着# l& p8 z* @$ R# G) N: \! _! e4 }2 z) `) j$ V$ x) m- z( V# D2 o$ G- ^( v8 o把头埋进臂弯7 o8 \+ k  J  j; j"" Y. g6 [  ~; d' C1 T7 ?/ x4 [5 T' g/ {/ I授奖词：| E) V"" ^% ]% H6 a4 u1 F9 G: j! s4 y; Y: Y"" H1 G8 `- m% Q1 A; e2 E在当下群星闪耀的年青一代女性写作者群落里 陆辉艳有决然不同的光芒和声音――它不是柔美的竖琴 而是金属的铜号。其新作《心中的灰熊》甚至具备了超越性别的坚硬、直接喝凌厉肌质。它沉静 冷峻 在小心翼翼的叙述里呈现细节化的真实 又曲折 回环 处处闪烁着超现实主义的光芒。有鉴于此 我们将第一届“青年文学•中国青年诗人奖”授予诗人陆辉艳女士。3 x3 K) v7 [9 Y# A6 u9 \/ P5 H: `5 Z  [5 o& y! i3 t' N: f* E' ?/ z# G| \6 K8 B/ l/ Z陆辉艳 广西作协会员 代表作有《静静伫立》、《缺席》等。* Y: E5 Q; n; ^# h  C7 k"" N( _$ h/ p& f7 w7 h( I| T9 C5 f- n  C- y"" m4 @6 D二、晴朗李寒《月光下的磨刀人》 2 C: I# C| ^' _'  * k- \| ~# ~# L8 W% m| ~| z! F+ O| L"" u9 L1 Y| I) ^* J. B7 P1$ g| r"" o| ]  u# a1 d6 W* ?' e7 ^: z% z: K* v! s0 r2 P% C0 e"" H7 o4 ^3 _8  1 d) x  J1 D我梦见 一个男人在月光下1 d  s- i8 s! r* S5 D. U| W& Y) P9 P2 w/ F: N$ C/ h4 z5 t' S' B"" X7 T磨着镰刀。+ R7 t* I- }/ u- d8 ?/ d8 A# f  i9 s1 Z4 E9 I: Q3 T+ `8 K5 {' M- t  ~8 m* @空空的院落被月光淹没 他低着头 2 e# a4 \' \  _. a% P4 u4 K( ]# W' @! {3 b8 V"" N0 {0 W; }; t* _(  ; d在磨刀石上刷啦刷啦地*  1 {# b% q| _* C* m' Z"" p( N6 k% q& ~( e; C; T5 d- r5 {) V. C磨着他的镰刀 他的身躯有节奏的摇曳 : b; L2 l2 f  R' b3 L' @| R| E; K' h' K: L$ u) h+ E: u8 _. N镰刀的锋刃 在石头上划出: B; a2 y: y  l# r6 u4 r2 e& p+ u5 K: T% i7 n: c6 C: v! q"" H1 O% e. n3 M: i- ^岁月的弧度。) V) F* u) b5 W* l: G9 K1 [6 j$ c% U- x' Y)  / Y  {2 R*  4 I. {  m8 i9 K% x$ @整个村庄的夜晚 除了偶尔的虫鸣 1 h7 h  H% p$ s2 w/ H0 T+ p. x4 Z"" j| x$ n$ B8 C3 r  b1 k! l( h6 p只响着他沙沙的磨镰声。( s4 B! M; c- M! C0 H* x( z/ n| Q9 X4 C9 t% a+ F7 w' C4 c- z: y0 k他 时而停下来 在石头上8 W/ G; S"" l1 O$ @* J8 N"" E6 i. U- P- w* Z"" w| k9 g) u8 a7 N! o洒一些水珠 时而用拇指轻轻试探一下; F"" B: \+ G8 V9 h' c! `+ f+ H| u& S| I! T$ j: D% E4 P/ P| v4 _' h锋刃+ d- ]7 ?4 D2 V1 q/ k3 t/ U* I9 `' N) y. F# H4 Q/ i8 {7 }) i% v) L"" }% o2 ^/ _. d$ b23 k"" I| w! [2 B' w- r3 s7 I5 i- T1 o% M1 a- k7  / j5 f1 r# O6 V) O( N| i月亮 也像一块光洁的磨刀石 6 J! f* ]! j9 y5 i8 e0 v$ s! _: a2 P1 q' _- e!  $ C9 y. @"" f-  - S% ~( }由圆满而渐渐残缺 它被谁的锋刃| V| U  V6 v6 n7 z' E1 d7 M1 O3 }  {3 D; T5 ?  X. W0 Q# ?| Q/ C越磨越单薄 越磨越弯 ! V% ^5 X4  - l5 G' j1 M. Z2 C3 b8 ~' b8 m3 r: R6 J& b5 X! P: }6 B# I3 N6 u  Q8 v; y"" ^最后 镰刀 磨刀石 月亮 这个男人$ x9 q4 }! Z& o7 W) `! R3 m) k% F/ H( y; H' q# Q8 w4 j8 N! L! P都有了相近的弧度。5 j& @| `6 }8 ]9 x+ G: i2 Y. P9 w  M$ l1 M/ D$ N+ Y+ K% m9 a3' }0 _) W. ~4 q6  8 O$ h1 ]# X9 x. v  ~0 e3 h* J  a& i$ }- {$ U. c9 M7 x这个男人 我不清楚他是谁3 d1 h' R+ v8 H: Z* ^"" B2 v5 S* C( K9 z. K. e3 q| G3 K8 a' _* T- [/ t  }. h也不知道 他将收割什么' U! w| z# O' c9 D% J4 x8 Y  r) ?% D/ C| v$ B) K4 K& _"" ~$ q! j3 G我只梦见 他坐在月光下( ?' J/ K7 s8 ]2 v+ e  q- a  u"" J8 k' W( w2 y"" I5 O. e一声不吭地磨着镰刀"" m3 V6 H. _  F! H: I0 w3 j| l3 l: j+ W+ _7 R# V- s| r2 Z"" E刷啦刷啦的声音在寂静的深夜| d- e) b; r2 `8 O"" c( N- m. e9 f# m0 V| V; b7 y6 `4 U+ A) @| e传出去很远很远% m! q2 n7 q) @4 C3 Q/ [. e- n) T  F3 j# ~3 D$ @7 E. U$ h2 j0  $ y0 \- f* L露水正集结到草叶上. l0 L. V3 p' s4  + E% E$ I8  - C& u$ R% B' V9 t4 G. E; S4 e/ T! \/ A* k( ^5 F0 }. `虫子的鸣叫也由浓渐稀# M$ E1 @9 w3 v"" y8 Z* I% B6 g  U7 ^  i) H% v+ z) w. ~( }$ u4 X+ Y5 U* k这个男人 还没有要停手的意思4 R9 Y# \"" Q; f  R4 ^/ h: m6 Y2 J* ^8 y( E| ~3 h( n7 @  u+ {4  我知道 他的镰刀已经很锋利了"" f! B2 k* i8 o# H! {- Q: N4 j% N1 f* w! A2 i# `  N& L0 H  Y% K# M"" T/ h' e4 Q' Y* E可是 他坐在月光下( ~' \2  2 h& s$ ?"" h( T2 u* t; M! V1 ]3 e5 \2 }2 l! d1 g/ n! F2 a佝偻着身子 倾注了全部的力气( l! d% Y6 f2 P1 p; `1 U& l  K$ Z3 o5 Y* ^  j( s* s% i- j' c* u8 ^& W( L8 c将一柄镰刀"" q0 ?5 t5 t) J9 A! a0 J& W8 M7 `0 p8 \5 u& N6 U: ~% [' M  u( Q2 V% D  T磨得越来越单薄( D  c% r2 I3 Y* S4 }8 ^) ]/ D8 C+ B0 J& I$ ^2 f  i2 W( i像秋风刮过树梢儿  l7 _3 r& Z! S4 R  L- B; ?/ ^* G3 O# r' l) }: x- s& L) q& E| W6 l9 H吹出清凉的寒意4 S8 D) q& k3 _7 y* @5  8 U; S/ _% y+ M"" V* k' ]0 N' y41 \0 ]* W! e3 Q% x+ _1 h$ n& \. N8 K| b8 g) R. T+ Z# T"" N  O; x2 f9 S2 P6 B月亮都隐没了 磨刀石也消损殆尽1 @! M"" c: }/ h# R  _) f5 k) r5 X: L5 W  m' J8 c: P- M' r) H1 j8 f9  ; v"" c黑色的楼群从四周包围上来 ' @"" j' A% r! w8 `! h% ~2 o: l1 o- `0 P# T1 z8 N% o5 i5 T已经没有庄稼可以收割了 * E0 W2 W9 i7 L3 k"" l$ o! P( J0 z: J9 k"" V0 _4 E0 y3 r) G"" O- ^; {这磨刀人的手中% t8 t4 w& u  Y4 M| \% L  Z% k7 P  P| ^"" d9 H6 Z4 J7 O$ ^& a$ g6 v& `7 b# l3 }也已经没有了镰刀 9 E5 P! e) D6 l| O+ F. C5 d% a* y( t8 I6 b; r| g) \' [  r# u5 s4 f; K  ?"" P他却仍旧向着虚空; D| @9 y. y5 D8 z6 D1 k; u3 A' Q/ `' @7 ^7 E$ A& ~* O! c8 w7 r. f做着磨刀的动作 他的嘴里发出( l"" U3 N3 f1 ?2 T( ~( Z"" k' \3 i# }5 @! X/ [$ q3 A$ F3 K- }/ u; ?"" f( Q8 a刷啦刷啦地 模仿着磨刀声。! K1 x5 F0 s+ j( C"" d( c4 J- r0 y| H8 k8 T  x  l) ^7 O* @) i( A: z; U此时 我才突然发现 + X: l6 x: c& R( q3 _4 [5 l- Q; w. H8 e+ E6 o# R5 K9 l# o$ s3 x6 c他的头 $ ?0 E5 j. N  \% x  O. p6 K; g) ^1 j8 z! u1 e# d& B$ L) L! V/ x3 v9 z已经白如小小的雪山。. p: w. ^: t! S/ w( O# D2 g"" h8 x# M* Y: o1 B' [$ j0 v| E8 L' T1 g# D/ [$ P  C( W授奖词：& z2 _6 d  `& O.  6 ?5 _! e! q* d0 j' C+ y4 ?8 F诗人晴朗李寒穷数载之功 呕心沥血 为中国读者奉献出了俄罗斯接触诗人阿赫玛托娃四卷本的诗歌全集 为中国当代诗歌写作提供了足可借鉴和学习的标杆 并将相同的尺度作用于自己的诗歌写作 写出了《月光下的磨刀人》这样的优秀之作 这些作品既保持了优美的抒情 又容身于当下现实 扎根于个人生活 表现出了诗人作为芸芸众生对生活的承受力和敏锐而广阔的精神世界 写出了个体生命不妥协的理想精神和独属于诗人的自我尊严。有鉴于此 我们将第一届“青年文学•中国青年诗人奖”授予诗人晴朗李寒先生。8 j6 y) @' _- j/  | l& ?5 {8 C2 M6 G8 H# A' c9 I1 ]: d2 h& c6 V9 b5 i0 T  _  l晴朗李寒 诗人 翻译家 河北省作协《诗选刊》杂志社编辑 代表作有《空寂与欢爱》等。' p& E1 @) t+ f6 z1 p( k$ N"" y( z  t1 J0 }5 g4 V"" X% F5 w# J* j& W. P+ P"" X) n; M三、黄明祥《从未有人走过》 9 M' l6 o- T| ^' D& k  \; E- {% [4 K* Q4 _9 l# b8 `6 S+ K7 q7 q; N# y我走过% L) _. I4 X"" e  f6 X# d6 C| u: e# S2 w. v/ k4 o"" Z:  . E0 v( O! t声音在脚底消失9 ]! F( `2 M- \1 x- s9 P: `  ~7 x; `0 z- n% c0 s! `/ @$ e6 x3 ?4 ~+ G; l8 K仿佛沉入水中# j7 A& [. q5 x2 p( o' F9 j2 F/ q. H1 a+ }& R9 `' ]% k  q4 v+ W* k8 z灰尘卷起小小的浪& g' j% e5 Q% b4 P9 i; U. s4  $ O% }. W| M% O6 D; }; w"" l7 K6 U7 ^; q- k# ?; u我忧心远行6 J; O$ H6 T$ d| y3 e$ r- f! b' n+ S1 q: L3 r  G9 K7 y! J$ i| [; u9 A; z0 _& K. i; J* M如果远行 浪会是一条河9 `9 F2 k4 g6 \$ y: }0 d: K) u  g( Y0 ?& L) B# v"" t流向海% T8 A( r& ^4 f( `$ n3 D/ Z0 s3 l. L8 r9 v9 J6 P5 Z$ \; V! O4 z9 t我害怕漂浮2 j; M& R) }3 ~"" w6 M% @/ E& R| T"" ^4  2 R) {4 M6 b' S2 P5 S不能寄望阳光成为灯塔' B6 L6 }% B; G- }3    y. L3 r1 S1 M- a- d6 h3 ]5 ^& e"" M5 O* Y| h将无边无际' @; b- o4 {& c| G1 }3 F1 d5 T& B( m- Z' W0 y! l4 E% H: c( _0 w3 P; Y: {照得毫无着落: N- p: x  u0 h3 M3 a$ d; f8 I3 G/ E' [( a. O1 C! \$ r/ N- m我只能漫步/ k: _+ F7 V9 x% J! F$ ]! g6  1 ]"" d& }  A; k- }: h4 q| V  C3 C7 _- C- E( y开一朵小花在走过的地方* V# f6 T0 O: m) G- U: P! h* v4 Q  x3 a4 f- r7 ]* J  I& m1 s3 D. U我驻足 等一棵树萌芽. n8 X  ~/ Y. Q! M( C| w$ i1 j( l6 t+ F1 ~| A| X0 }0 w2 g走过的地方) o8 ?  I/ D# F| N+ T- @  {' \+ ?) ]9 F| j# k: J# [- U- o5 C6 \$ T# r5 d! e. y9 I走着走着就走成了荒原( V9 X6 h3 y( Y* K9 u| c* T"" ^0 y2 P"" j4  * z0 `) }! L' U  ?5 J7 ~- x下一片连上上一片+ M# u4 I% v( S( Z: f; }8 U7 M7 R( x. e: F# p- J% x9 U6 I0 M9 K年轻的事物都在老去. H$ `) \5 T2 J1 e3 ]$ V  l1 ^$ ]4 V9 x  `# H  G) U; m$ I6 m2 E老去的 在想走前的事| _' B) l| o0 M: N4 B' m+ J1 v7 }# Q/ C; k# W5 B# M# U7 S) i3 d  s2 f3 Y& H2 I8 d| w仿佛从未有人走过+ R5 P& V: [( V1 e. t8 A& @! f' [: R% u9 N& k  f: E1 V9 T8 a3 A) o! B9 P: Q# D* @% e4 v8 u授奖词：; H2 w0 g| f) v) V; n! _2 S0 J+ R) ~5 ^- j; \# O5 ?# I7 a* c$ a) v! G"" \- G9 U  J诗人黄明祥在自己并不长久的诗歌写作生涯里 从一开始就表现出了独特的个性和勇气。其组诗《从未有人走过》简约、淡远而又深情、内敛 他专注地使用着自己独特的语言谱系 他的专注里有着窥伺者的犀利和精准 并坚持指向事物内部的秘密。这秘密当然不是故事本身 而是对世界的发现和再造 以及对自我“何来何去”的形而上思考。有鉴于此 我们将第一届“青年文学•中国青年诗人奖”授予诗人黄明祥先生。4 X# ^# L  T$ d& t. ~/ K/ j2 W' X' d' ?8 l9 L( P7 V2 i5 J+ }黄明祥 诗人 收藏家、艺术评论人 《十月》杂志艺术主持人 代表作有《中田村》、《铁匠》等。. J; I8 f  [0 ?3 E/ }) z# n3 y"" c  ^| t  C  c  j* E书记处书记| 社会实践| 湖南湘西| 吉狄马加| 南国早报"|http://www.ngzb.com.cn/forum.php?mod=viewthread&tid=1251339&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline|2015-10-31
其他媒体|2096464174|zhidao_baidu|电脑/网络 > 笔记本电脑|ZHO|2015-11-03 01:18:01|"东风雪铁龙世嘉1|6l品尚型和起亚k3标配|那个更优秀"|来自：手机知道汽车|http://zhidao.baidu.com/question/1896179845711881780.html?fr=qlquick&entry=qb_list_default|2015-11-03
其他媒体|2128220164|hexun|水煮爱车|ZHO|2015-11-20 18:17:02|哈弗H6改装TEC和ARC音响――武汉歌德|　　旅行 在意的不是沿途的风景 风景太多 我们无法一一记起 我们在意的是徜徉在风景之中的心情和留恋。音乐 在意的不是它的出处 旋律太多 我们无法一一感受 我们在意的是它给予我们心灵的那一份慰藉与感动。一套好系统的升级 在给予自己内心最大欢愉的同时 也给社会带来不少的正能量。下面我们就一起来欣赏一下武汉歌德带来的这套充满正能量的发烧系统吧！首先我们来看一下升级配置：替换原车主机 改用阿尔派9887 外加一台阿尔派H800处理器来稳定音源 前声场升级意大利TEC SQ6/K3三分频 后声场升级TEC SQ6/K两分频 一只低音辅助声场 驱动则由三台美国ARC旗下具有“黑匣子”之称的KS系列来担任 光看配置 就能感受到它能量的波动 如此发烧级的升级套装 最后到底会为我们呈现出一场怎样的音乐盛宴呢！小编我也不得而知 想要知道答案 就请大家跟随我一起来探索一下吧！　　　　哈弗H6汽车音响升级 全面改装TEC和ARC音响　　　　前声场意大利TEC SQ6/K3高中音单元A柱倒模安装效果　　　　前声场意大利TEC SQ6/K3中低音单元安装效果　　　　中控台纵览　　　　后尾箱安装整体效果　　　　阿尔派H800信号处理器安装效果　　　　美国ARC功放 KS1500.1安装完成效果图　　　　尾箱器材安装排布井井有条 在加上在七彩变幻灯光的映照下 使得尾箱更是颇具几分神秘色彩。　　　　系统点评：当最后一道工序调音落下帷幕 昭示着H6音响升级的过程已全部完成 也可以说是TEC与ARC金牌组合又一发烧系统新鲜出炉 店家专业的改装技术与严谨的工作态度让人无可挑剔 完美的SQ音 再有“黑匣子”之称的KS系列功放的驱动下 其音质的发挥更显得如鱼得水 就好比是伯乐遇上了千里马 两者惺惺相惜 事半功倍 轻松为车主共同谱写一段新的音乐传奇。　　 　　哈弗H6音响改装配置：　　主  机：阿尔派9887　　处理器：阿尔派H800　　前声场：意大利TEC SQ6/k3三分频　　后声场：意大利TEC SQ6/K两分频　　超低音：K牌L5　　功放一：美国ARC KS300.4四路功放　　功放二：美国ARC  KS300.2两路功放　　功放三：美国ARC KS2500.1单路超低音功放　　线  材：霸克2号电源线 佰利2M音频线 霸克喇叭线查看更多精彩内容请进论坛首页|http://bbs.hexun.com/post_111_9033141_1_d.html|2015-11-20
其他媒体|2128628849|zhidao_baidu|电脑/网络 > 硬件 > 内存|ZHO|2015-11-20 22:46:03|东风悦达起亚k3有没有前后防撞钢梁有的话防撞钢梁的厚度是多少|来自：手机知道生活东风悦达起亚k3有没有前后防撞钢梁有的话防撞钢梁的厚度是多少|http://zhidao.baidu.com/question/490855599336517772.html?fr=qlquick&entry=qb_list_default|2015-11-20
其他媒体|2227075063|zhidao_baidu|生活 > 购物|ZHO|2016-01-17 17:07:15|起亚k3飞歌g6s导航怎么和手机互联|赛车|http://zhidao.baidu.com/question/427521547981401772.html?fr=qlquick&entry=qb_list_default|2016-01-17
其他媒体|2227403820|zhidao_baidu|电脑/网络 > 硬件 > 硬盘|ZHO|2016-01-17 21:27:14|起亚k3怎么锁了会自动四灯全闪门也会开|汽车我是东风悦达起亚k3车怎么锁了会自动四灯全闪门也会开。|http://zhidao.baidu.com/question/555265431109026052.html?fr=qlquick&entry=qb_list_default|2016-01-17
其他媒体|2320021562|bitauto|易车 > 问答 > 问题分类|ZHO|2016-03-09 09:10:01|是北京现代朗动好还是起亚k3好|是北京现代朗动好还是起亚k3好     提问者：汽车报价大全**********  分类：  现代  朗动  其他  浏览[8] 来自：易车手机客户端  2016-03-09 08:04  举报   是北京现代朗动好还是起亚k3好|http://ask.bitauto.com/detail/6279806/|2016-03-09
其他媒体|2320151350|zhidao_baidu|电脑/网络|ZHO|2016-03-09 10:40:01|东风悦达起亚k3手动挡多少钱sohu|汽车|http://zhidao.baidu.com/question/1433505116115937139.html?fr=qlquick&entry=qb_list_default|2016-03-09
其他媒体|2321111074|bitauto|易车 > 问答 > 问题分类|ZHO|2016-03-09 20:14:02|东风悦达起亚k3手动挡多少钱sohu|东风悦达起亚k3手动挡多少钱sohu     提问者：易车网友 分类：  东风  买车  报价  浏览[2]  2016-03-09 19:12  举报|http://ask.bitauto.com/detail/6282375/|2016-03-09
其他媒体|2349149996|zhidao_baidu|电脑/网络 > 硬件 > 硬盘|ZHO|2016-03-25 10:05:01|东风悦达起亚k3s怎样装车牌视频|汽车|http://zhidao.baidu.com/question/563054935698418324.html?fr=qlquick&entry=qb_list_default|2016-03-25
各大媒体|2349415329|enorth|汽车频道|ZHO|2016-03-25 12:59:01|悦达起亚k3现车优惠4万 国产口碑韩系轿|　　【网上车市天津滨海行情.原创】近日获悉 东风悦达起亚k3现车到店发售中 国产紧凑型轿车全系优惠4万最新独家促销价格。东风悦达起亚k3配置丰富手续齐全 具体颜色和配置请致电商家咨询 一手贸易商拒绝中间加价 更多优惠尽在北京诚远诚丰汽车销售公司 如您对本车感兴趣 欢迎致电咨询 购车热线：　　***********刘经理　　具体车型以及价格如下：　　本车报价：　　外观方面 东风悦达起亚k3在前脸的设计上十分突出力量感和线条的精炼 采用起亚旗舰车型K9的镀铬直瀑式竖条进气格栅 视觉感受更为大气、稳健 后尾组合尾灯和外后视镜集成转向灯都采用LED设计 再配合LED日间行车灯 彰显出浓厚的科技感以及时代感。　　细节方面 东风悦达起亚k3的超长轴距更打造出同级别最大乘用空间 充分保障了驾乘舒适性。K3还配备了电动通风真皮座椅、双区恒温空调、一键启动、高级音响系统等同级罕见的科技 充分体现出K3配置的丰富和越级。　　内饰方面 东风悦达起亚K3简约内饰 完满组合时尚先锋梦之队。K3内饰做工精致 真皮座椅、方向盘、门护板、仪表盘等皮质包裹 触感细腻高贵 工艺超越同级。K3的配置套餐也极具智能感 与K3族群“科技控”的前瞻审美观无缝衔接。　　配置方面 东风悦达起亚k3还搭载了起亚最新的1.6L伽马D-CVVT和1.8L Nu D-CVVT两款发动机 最大功率分别达到128马力和146马力 动力强劲且燃油经济性突出。配合先进的6速手自一体变速箱 操控随心 能很好的开发车主驾驭热情。【网上车市天津滨海行情.原创】　　更多详情请点击： http://binhai.cheshi.com/网上车市滨海车市　　温馨提示：以上购车优惠信息由天津滨海综合经销商提供 仅供购车参考；由于行情因素价格浮动较大 具体车辆成交价格请致电商家获取最新报价；优惠行情可查阅网上车市天津滨海经销商报价后台 告知对方信息来源于网上车市将有更多优惠。|http://auto.enorth.com.cn/system/2016/03/25/030886245.shtml|2016-03-25
其他媒体|2350225543|bitauto|易车 > 问答 > 问题分类|ZHO|2016-03-25 22:14:01|东风悦达起亚k3s怎样装车牌视频|东风悦达起亚k3s怎样装车牌视频     提问者：易车网友 分类：  东风  其他  浏览[3]  2016-03-25 21:12  举报|http://ask.bitauto.com/detail/6345539/|2016-03-25
기타|2416104604|Autohome review|혼다 어코드(雅阁)|ZHO|2016-05-01 00:24:12|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=111&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-01
기타|2416273106|Autohome review|혼다 어코드(雅阁)|ZHO|2016-05-01 03:03:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=112&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-01
기타|2416597534|Autohome review|혼다 어코드(雅阁)|ZHO|2016-05-01 10:53:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=113&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-01
기타|2416759558|Autohome review|혼다 어코드(雅阁)|ZHO|2016-05-01 13:05:03|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=114&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-01
其他媒体|2416800057|bitauto|易车 > 问答 > 问题分类|ZHO|2016-05-01 13:39:03|东风悦达起亚k3。 1.6l自动顶配10.88。 怎么样。同|东风悦达起亚k3。 1.6l自动顶配10.88。 怎么样。同     提问者：汽车报价大全**********  分类：  买车  选车  浏览[9] 来自：汽车报价大全  2016-05-01 12:25  举报   东风悦达起亚k3。 1.6l自动顶配10.88。 怎么样。同等价位还能考虑什么。 地址是在黑龙江。|http://ask.bitauto.com/detail/6499506/|2016-05-01
기타|2417074998|ngzb|新闻互动|ZHO|2016-05-01 17:14:02|柳州：创作山歌MV 民警爆红网络|"马上注册 结交更多好友 享用更多功能 让你轻松玩转南宁您需要 登录 才可以下载或查看 没有帐号？立即注册  x创作山歌MV 民警爆红网络主要宣传各种法律法规 网友点赞“太有才”南国早报网―南国早报记者 陈新援3 e9 i& {  T1 g& i# D'  155.jpg (125.4 KB| 下载次数: 8)下载附件 保存到相册1 小时前 上传韦茂个人原创山歌《山歌唱起枪弹炮》的视频截图。0 c. \+ t# W"" ]) n* }　　最近一部名为《山歌唱起枪弹炮》的视频“刷爆”了柳州市民的朋友圈 这首歌以宣传缉枪制爆为主要内容 看似严肃的主题 被用桂柳话山歌唱出后 竟然令无数人着了迷 短短两天 点击量就超过了10万 好评如潮。那么 这究竟是一首什么样的歌 唱山歌的人是谁？这首歌又是怎样创作出来的呢？) ^8 N5 o2 }0 n/ w( J5 M: ~0 s& C& N; ?"" ?4 D; h　　幽默山歌获点赞& n| O* ^7 R  x6 Z* i% ?0 d3 z2 q/ @/ N+ W$ w( P/ E9 v"" X　　“这个老派（警察）唱的山歌真有趣 太有才了！”最近 在柳州市民的朋友圈里 不少人都在竞相转发一则视频。视频中 一名身穿警服的男子 一边弹奏电子琴  一边摇摆着唱起山歌。8 Z"" I& F4 q) P' c5 V! _& F"" k3 [5 p"" h! v0 x9 O　　“乱玩枪弹更可怕 3 Y2 ~$ a0 Y4 X| v$ y2 O. N; F# I3 ^7 I* w% x# y! t( Z$ ^　　惹出麻烦你头大。1 t( _- p- R) X4 a1 W: v% v& S4 a"" A/ A( R* ^　　子弹铁砂没长眼（哩） | Z1 b5 A3 Q. z) k# p7 b% u"" ]"" m/ H) G0 D0 I　　伤人毁物几鬼险。)  # F( H& ?$ X* s9 k( n/ H8 h'  1 I7 @7 m3 S2 u3 O/ K2 O| t) E　　你自己看（勒）你自己看（勒）你克玩这种 % @1 I"" {( }6 _% ?+ b; z& D* R1 w( L% t  V( g　　误伤自己你倒霉（呀） )  7 _4 s$ U- R  e- g8 ?7 T* Q6 N  J1 j6 ~* {% H7 `　　打到别人要命赔。9 l. t- J1 E4 e6 X$ e1 b6 U: H# @' P"" w7 V4 ~　　要是藏有枪和弹哩 . f"" M9 i9 i# F* c-  $ o6 C( y2 g  O; K$ ~　　害人害己屁股宽。8 P4 q+ `/ Y: X' ]! t1 o5 t) {* K. m/ k- x4 j　　白：（哎呀）我见（哩）屁股宽过大海（哩哦）”。/ ?1 P9 A! ?% ~% r2 j"" L% c* A3 a' {9 ]　　桂柳话唱腔 配合着诙谐幽默的旁白 听罢令人忍俊不禁。一名网友评价：如此宣传没有生硬刻板的说教 形式活泼 语言朴实又不乏幽默 非常接地气 让人在会心一笑的同时 也在脑海里记住了宣传的内容 是创新之举 点赞！. s$ u8 l! L6 C# M+ a( `; Q| \4  9 H; ?: _# U& }　　还有网友评价 这首歌初听起来觉得有点“土” 不过细细听完 觉得很有意思 后来竟着魔般反复听了好几遍。记者看到 这首MV被某微信公众号转载后 在短短两天时间 点击量已经超过10万 点赞近千。6 ^! l/ Z7 y| h- d  @/ Q: u6 o! l( t; ^. Q# B& `　　用业余时间录制* J- B7 q; X# N% S8 y0 r| j% w( e5 g7 M　　据了解 这首MV的创作者和表演者 是柳江县公安局指挥中心教导员韦茂。韦茂从事公安宣传工作多年 2012年开始通过壮语歌曲向群众宣传法律、宣传公安工作 受到当地百姓追捧 被当地群众称为“警察歌星”、“壮乡民警歌星”。  A6 W- r-  / ^  p: x5 X6 ]7 ?"" m"" d# {0 F/ g5 J2 K0 H"" ~　　“都是业余时间制作的。”4月30日 韦茂在接受采访时说 这首歌其实这是一首“老歌”。2015年10月13日起 公安机关缉枪制爆“神剑1号”专项行动在广西各地开展 从事宣传工作的他 也开始思考采用什么新方式进行相关宣传。山歌是少数民族地区群众喜闻乐见的一种艺术形式 于是他决定把相关的法律和政策融入山歌中来宣传。从构思、谱曲、写词到录制、混响、后期剪辑 几易其稿 反复修改 前后先后花了一个多月时间 全由他一人搞定。( a% e| M. S) m5 l% w( ~. M# V5 Z6 M; B* S9 O! J　　韦茂说 这则视频拍摄地点在他家里 弹奏用的电子琴是他女儿“淘汰”的 背景就是他家的一面白墙壁。没有华丽的舞台 也没有讲究的灯光布景和音效 一切都是“原生态”。- x- r  e1 y3 }7 Y"" ^% v( I: x4 {: A* F1 b　　他首先用录音设备将歌曲和音乐录下来 通过电脑制作好歌曲 然后 再在房间内架起电子琴和摄像机 戴起耳麦 和着音乐 一边弹唱一边“自拍”。"" o6 H0 e/ c6 A' X( I"" [' Y4 r5 u/ n$ f| f# N5 E1 T1 c0 D' K　　“反复录制了好几遍才成功。”韦茂说 由于是原创的歌曲新歌 要一次拍摄成功非常困难。就这首歌 他反复弹唱录制了好几遍 并且在后期电脑制作时花了比较大的功夫才最终制作完成。; A1  % H3 t: Y5 ?7 n/ m4 ?"" ~' O! {| s7 I% U( N5 N"" b9 G( Z4 P( U; N　　2015年11月底 韦茂将制作好的MV上传到了土豆网 一下就有近3万的点击量 好评如潮。最近 有人将他的视频上传到了腾讯视频上 并在朋友圈中进行了转载 结果再次爆红。# J- ^. c3 i5 W) K/  "" V- B; l& p; B9 Y　　歌曲成“盗版”热门) C9  * G1 k9 M"" }( _- y* K2 f* f) I0 Y8 H　　其实 这个已不是韦茂第一次制作这类宣传视频 早在2014年 他创作的一首奉劝群众远离毒品的《禁毒壮语歌》一度风靡网络 短短几天时间 点击量就超过7万。柳江县禁毒办和柳江县电视台得知后 立即给予大力支持 他们派出专业人员为韦茂录制了MV。这首MV于当年“6・26”国际禁毒日当天在县人民广场首发时 就引来近千名群众的围观。7 K  Y! x( _0 B4 l7 h6 `; H) ?| G4 V% j　　韦茂创作的歌曲蕴含着浓郁的乡土气息 语言朴实、形式活泼 内容浅显易懂 非常受欢迎 他的“粉丝”已遍布全国各地 在柳江县更是拥有大量忠实的“粉丝” 不少人还专门找韦茂讨要歌碟 韦都热情奉送。韦茂说 到目前 他已送出上千张光碟 光刻录机都刻坏了几台。$ L! s6 j"" K2 H$ `# L) J8 }2 Q4 l9 j8 k; G) h& x  b3 e　　为了让更多人听到他的歌 他在土豆网上注册了名为“琴心画意”的账号 专门用于发布他的原创歌曲。2 i) w! E# ~- b7 `6 ^) R6 }- @; I| R& x| V8 Q4 Z' L　　现在 韦茂已经创作了二三十首用壮语和桂柳话弹唱的歌曲 这些歌曲中 有劝导群众远离“六合彩”的 有宣传公安工作的 也有祝福美好生活的。最新的一首是今年3月份创作完成的《家安天网人财安》 目前该视频在土豆网上点击已近万。1  3 p5 e0  + n* P: D  ~% v# X/ u4 P8 I3 L　　一些小商贩也嗅到了“商机” 从网上下载韦茂的歌曲 刻成光碟在县城里销售 结果非常抢手。一般的光碟 10元钱3张 而韦茂的歌曲光碟10元两张。  ]# e# s7 g| B8 F  ?% P# f: d# A/ _$ B4 Z)  ) V  V& f　　虽然自己创作的歌曲被盗版 可是韦茂并不打算深究。他说 创作这些歌曲的目的就是为了宣传相关的法律法规 能让更多的人听到这些歌 通过歌曲学法、懂法、用法 这也是好事。( Y"" I0 K- U3 y7 q1 U. k+ X"" L7 V* N0 j% r% _% b; S0 l! O南国早报| 电子琴| 主题| 朋友| 柳州"|http://www.ngzb.com.cn/forum.php?mod=viewthread&tid=1284524&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline|2016-05-01
其他媒体|2420099721|cqsb_cqnews|华龙网新闻中心-国内频道|ZHO|2016-05-03 10:41:07|与兰州舰一起演练的这些外国舰艇实力如何？(图)|5月1日 参加东盟防长扩大会议海上安全与反恐联合演习-2016的中国海军南海舰队兰州舰抵达文莱穆阿拉港 此前已有五艘参演舰艇抵达 分别是美国海军DDG-63斯特西姆号、俄罗斯海军572维诺格拉多夫海军上将号、韩国海军981崔莹号、印度海军L24埃拉瓦特号和越南海军HQ381号巡逻艇。本次各国派遣来参与联演的舰艇中 有中美新锐的“盾舰”两艘 俄罗斯大型反潜驱逐舰一艘 韩国通用驱逐舰一艘 印度登陆舰一艘以及越南海军巡逻艇一艘。其中 DDG-63“斯特西姆”号服役于美国海军第七舰队第15驱逐舰中队 属美国海军主力驱逐舰“阿利伯克”级FlightⅠA型 为伯克级早期型号 最初作为提康德罗加级巡洋舰的低成本高效能版存在 是美国海军第二级搭载宙斯盾系统的防空舰。全舰主要以宙斯盾系统为核心 武备方面主要有十二组共96单元Mk41垂直发射系统 一门Mk45127mm舰炮 两座四联装鱼叉导弹发射架 两座Mk32三联装324mm鱼雷发射器以及两座密集阵近防系统。作为美军主力驱逐舰 伯克级功能全面 作战能力强大。对空方面“标准”舰空导弹配合“密集阵”近防系统组成两层防空网 对海则有“鱼叉”反舰及“阿斯洛克”反潜导弹 Mk32鱼雷发射管发射的Mk46轻型反潜鱼雷 对陆攻击则有“战术战斧”远程陆攻巡航弹为主力 以及Mk45127mm炮作为对陆、对海攻击的补充。可以看出 伯克级作为美国海军90年代的“新生代” 是现今以及未来相当一段时间内的舰队主力 各方面性能均衡而强大 尤以防空和对陆攻击能力较为突出 其先进的宙斯盾系统和远程的战斧导弹提供了远超其他国家普通驱逐舰的强大作战能力。FlightⅠA型由于没有机库 反潜能力相比后期型号稍弱 在战斧反舰型号相继被取消以及LRASM未服役的情况下 本舰对水面舰攻击能力也只是一般水平。但综合来看 仍然是本次联演中战斗力最为强大的舰艇之一。【1】【2】【3】【4】【5】下一页|http://news.cqnews.net/html/2016-05/03/content_36819341.htm|2016-05-03
기타|2420099788|ifeng_news|凤凰网资讯 > 滚动新闻|ZHO|2016-05-03 10:41:07|与兰州舰一起演练的这些外国舰艇实力如何？|原标题：与兰州舰一起演练的这些外国舰艇实力如何？东盟身旁的大国舰影——参加东盟防长扩大会议海上安全与反恐联合演习-2016的舰艇解析■国防科技大学国际问题研究中心 青晨 李佑任5月1日 参加东盟防长扩大会议海上安全与反恐联合演习-2016的中国海军南海舰队兰州舰抵达文莱穆阿拉港 此前已有五艘参演舰艇抵达 分别是美国海军DDG-63斯特西姆号、俄罗斯海军572维诺格拉多夫海军上将号、韩国海军981崔莹号、印度海军L24埃拉瓦特号和越南海军HQ381号巡逻艇。本次各国派遣来参与联演的舰艇中 有中美新锐的“盾舰”两艘 俄罗斯大型反潜驱逐舰一艘 韩国通用驱逐舰一艘 印度登陆舰一艘以及越南海军巡逻艇一艘。其中 DDG-63“斯特西姆”号服役于美国海军第七舰队第15驱逐舰中队 属美国海军主力驱逐舰“阿利 伯克”级FlightⅠA型 为伯克级早期型号 最初作为提康德罗加级巡洋舰的低成本高效能版存在 是美国海军第二级搭载宙斯盾系统的防空舰。全舰主要以宙斯盾系统为核心 武备方面主要有十二组共96单元Mk41垂直发射系统 一门Mk45 127mm舰炮 两座四联装鱼叉导弹发射架 两座Mk32三联装324mm鱼雷发射器以及两座密集阵近防系统。作为美军主力驱逐舰 伯克级功能全面 作战能力强大。对空方面“标准”舰空导弹配合“密集阵”近防系统组成两层防空网 对海则有“鱼叉”反舰及“阿斯洛克”反潜导弹 Mk32鱼雷发射管发射的Mk46轻型反潜鱼雷 对陆攻击则有“战术战斧”远程陆攻巡航弹为主力 以及Mk45 127mm炮作为对陆、对海攻击的补充。可以看出 伯克级作为美国海军90年代的“新生代” 是现今以及未来相当一段时间内的舰队主力 各方面性能均衡而强大 尤以防空和对陆攻击能力较为突出 其先进的宙斯盾系统和远程的战斧导弹提供了远超其他国家普通驱逐舰的强大作战能力。FlightⅠA型由于没有机库 反潜能力相比后期型号稍弱 在战斧反舰型号相继被取消以及LRASM未服役的情况下 本舰对水面舰攻击能力也只是一般水平。但综合来看 仍然是本次联演中战斗力最为强大的舰艇之一。|http://news.ifeng.com/a/20160503/48661306_0.shtml|2016-05-03
기타|2420317514|southcn_news|中国|ZHO|2016-05-03 12:47:12|与兰州舰一起演练的这些外国舰艇实力如何？|　　东盟身旁的大国舰影　　——参加东盟防长扩大会议海上安全与反恐联合演习-2016的舰艇解析　　■国防科技大学国际问题研究中心 青晨 李佑任　　5月1日 参加东盟防长扩大会议海上安全与反恐联合演习-2016的中国海军南海舰队兰州舰抵达文莱穆阿拉港 此前已有五艘参演舰艇抵达 分别是美国海军DDG-63斯特西姆号、俄罗斯海军572维诺格拉多夫海军上将号、韩国海军981崔莹号、印度海军L24埃拉瓦特号和越南海军HQ381号巡逻艇。　　本次各国派遣来参与联演的舰艇中 有中美新锐的“盾舰”两艘 俄罗斯大型反潜驱逐舰一艘 韩国通用驱逐舰一艘 印度登陆舰一艘以及越南海军巡逻艇一艘。　　其中 DDG-63“斯特西姆”号服役于美国海军第七舰队第15驱逐舰中队 属美国海军主力驱逐舰“阿利伯克”级FlightⅠA型 为伯克级早期型号 最初作为提康德罗加级巡洋舰的低成本高效能版存在 是美国海军第二级搭载宙斯盾系统的防空舰。全舰主要以宙斯盾系统为核心 武备方面主要有十二组共96单元Mk41垂直发射系统 一门Mk45 127mm舰炮 两座四联装鱼叉导弹发射架 两座Mk32三联装324mm鱼雷发射器以及两座密集阵近防系统。作为美军主力驱逐舰 伯克级功能全面 作战能力强大。对空方面“标准”舰空导弹配合“密集阵”近防系统组成两层防空网 对海则有“鱼叉”反舰及“阿斯洛克”反潜导弹 Mk32鱼雷发射管发射的Mk46轻型反潜鱼雷 对陆攻击则有“战术战斧”远程陆攻巡航弹为主力 以及Mk45 127mm炮作为对陆、对海攻击的补充。　　可以看出 伯克级作为美国海军90年代的“新生代” 是现今以及未来相当一段时间内的舰队主力 各方面性能均衡而强大 尤以防空和对陆攻击能力较为突出 其先进的宙斯盾系统和远程的战斧导弹提供了远超其他国家普通驱逐舰的强大作战能力。FlightⅠA型由于没有机库 反潜能力相比后期型号稍弱 在战斧反舰型号相继被取消以及LRASM未服役的情况下 本舰对水面舰攻击能力也只是一般水平。但综合来看 仍然是本次联演中战斗力最为强大的舰艇之一。|http://news.southcn.com/fu/content/2016-05/03/content_147027997.htm|2016-05-03
기타|2434298109|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-11 00:01:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=20&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-11
기타|2434510644|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-11 02:32:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=21&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-11
기타|2434573312|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-11 03:41:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=167&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-11
기타|2434573352|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-11 03:41:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=12&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-11
기타|2434854076|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-11 09:24:02|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=168&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-11
기타|2434891953|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-11 09:53:03|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=13&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-11
기타|2435045708|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-11 11:25:09|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=22&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-11
기타|2435662681|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-11 17:11:02|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=169&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-11
기타|2435663196|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-11 17:11:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=14&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-11
기타|2435727072|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-11 17:44:04|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=170&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-11
기타|2435790616|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-11 18:16:05|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=15&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-11
기타|2436205291|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-11 22:11:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=32&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-11
기타|2436313078|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-11 23:14:02|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=171&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-11
기타|2436313343|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-11 23:14:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=16&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-11
기타|2436367122|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-11 23:47:15|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=172&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-11
기타|2436367419|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-11 23:47:16|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=17&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-11
기타|2436368364|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-11 23:47:17|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=34&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-11
기타|2442042307|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-15 00:15:04|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=10&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-15
기타|2442075778|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-15 00:42:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=41&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-15
기타|2442112027|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-15 01:14:02|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=12&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-15
기타|2442176489|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-15 02:15:01|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=13&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-15
기타|2442251586|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-15 03:55:01|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=88&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-15
기타|2442514633|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-15 10:41:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=187&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-15
기타|2442515000|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-15 10:41:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=32&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-15
기타|2442641978|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-15 12:27:59|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=89&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-15
기타|2442655506|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-15 12:39:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=188&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-15
기타|2442655918|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-15 12:39:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=33&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-15
기타|2442937000|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-15 16:20:02|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=90&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-15
기타|2442971520|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-15 16:45:02|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=14&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-15
기타|2443076322|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-15 17:58:01|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=91&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-15
기타|2443124556|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-15 18:31:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=42&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-15
기타|2443228794|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-15 19:49:01|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=15&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-15
기타|2443412927|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-15 22:09:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=44&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-15
기타|2443434219|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-15 22:25:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=53&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-15
기타|2443439555|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-15 22:28:02|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=16&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-15
기타|2443463384|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-15 22:46:02|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=92&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-15
기타|2443467332|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-15 22:49:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=189&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-15
기타|2443467702|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-15 22:49:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=34&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-15
其他媒体|2443475820|zhidao_baidu|生活 > 生活常识|ZHO|2016-05-15 22:55:02|东风悦达起亚k3最低配裸车多少钱|汽车|http://zhidao.baidu.com/question/1821390504309690108.html?fr=qlquick&entry=qb_list_default|2016-05-15
기타|2443485127|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-15 23:02:01|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=8&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-15
기타|2443526307|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-15 23:34:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=54&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-15
기타|2443526404|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-15 23:34:01|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=9&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-15
기타|2443543930|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-15 23:47:36|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=93&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-15
기타|2443558183|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-15 23:58:01|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=17&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-15
기타|2456879471|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-23 00:53:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=216&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-23
기타|2456879876|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-23 00:53:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=65&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
其他媒体|2457093023|chinatimes|財經 RSS|ZHO|2016-05-23 05:23:02|銀行圈粉 展開大作戰|"國銀「圈粉」時代來臨。進入Bank3.0後 銀行從過去搶財管客戶 轉向搶社群鄉民 「圈粉」大戰已然開打。目前圈粉最積極者 莫過於中信銀、國泰世華銀、花旗銀和永豐銀 各家除了力拚臉書人氣 也大舉經營網路社群 就是要鎖定更多年輕客層。有別於過去的自營粉絲團 圈粉指的是直接和現存粉絲團合作 把粉絲團的粉絲變成銀行客戶。像是中信銀就與GOMAJI還有iCHEF合作「圈」美食族、與EZTABLE點「圈」禮券族、與Pi行動錢包合作「圈」社群電子商務族。  中信銀消金主管指出 以GOMAJI為例 透過「夠麻吉卡APP」以信用卡付款 消費者不需更換手機 只要憑QR Code掃描即可完成信用卡支付 讓GOMAJI的客戶都可使用中信卡。永豐銀第三方支付平台「豐掌櫃」時則與PIXNET合作 推動社群商務 PIXNET DIGITAL MEDIA旗下龐大的痞客邦會員可直接安裝豐掌櫃APP在部落格中 讓永豐銀的代收代付服務立刻滲透到社群手機。國泰世華銀則與社群工具LINE Pay合作 提供購物金；並在Yahoo、PChome、淘寶網等購物商城提供特殊折扣或回饋金 並在臉書與臉友互動 啟動「大圈粉」行動。花旗銀行則是祭出「揪團刷卡」搶優惠 最令卡友瘋狂的是「月月可抽BMW X3系列休旅車」 活動推出僅20天就超過6|000團的花旗好友圈被建立 短短4個月內揪出18|000團 最大團超過9|000人。(工商時報)    關鍵字：臉書"|http://www.chinatimes.com/newspapers/20160523000087-260205|2016-05-23
기타|2457283284|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 09:38:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=112&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2457283478|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 09:38:04|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=42&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-23
기타|2457370483|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 10:40:03|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=113&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2457370705|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 10:40:03|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=43&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-23
기타|2457443089|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-23 11:26:02|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=121&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-23
其他媒体|2457456650|zhidao_baidu|电脑/网络|ZHO|2016-05-23 11:33:02|东风悦达起亚k3汽车15款和16款配置有什么区别|汽车|http://zhidao.baidu.com/question/811720771469320812.html?fr=qlquick&entry=qb_list_default|2016-05-23
기타|2457543447|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-23 12:24:16|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=123&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-23
기타|2457612724|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 13:07:19|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=115&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2457612938|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 13:07:19|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=45&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-23
기타|2457670335|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-23 13:44:02|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=125&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-23
기타|2457675759|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-23 13:48:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=217&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-23
기타|2457675938|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-23 13:48:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=66&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
各大媒体|2457686647|qc188|车主说车 > 紧凑型车|ZHO|2016-05-23 13:55:02|早已下定决心 谈现代领动1.6L提车心得|"话说从19号到今天也快一周了 碰巧今天25号（农历3月19）是我跟老婆结婚4周年 晚上的好好庆祝庆祝！写到这里不知从何写起了！先说说有购车计划到购车这段辛苦流程吧 15年春节老丈人一家来杭州过年 说起谁谁谁又买车了！现在孩子到杭州读书出去玩一家没车也不方便！我夫人就说现在滴滴优布打车这么便宜又方便 说到滴滴优布我想想自己上班休息时间这么多（白夜休休 基本上上一个白班休息3天 夜班就是睡觉）！最后和老婆商量没事可以跑跑滴滴或优步 想想自己拿驾照一年半了都没有摸过车 30岁的男人了现在没车以后肯定会有的 早买早享受吧 这之后就有了购车计划 预算在13万左右。问了身边同事买什么车好 都说的五花八门?? 有一个同事直接告诉我买车买自己喜欢的 问别人问不出来的！你买50w车都会有人说不好！出门天天看到楼下房东这辆索8 老婆也感觉这车线条不错 挺漂亮的（对车不怎么懂 只能先看外观了） 上百度一搜价格超出预算 于是天天在小区里转悠看看有没有什么好看的车！首先说明本人暂不考虑日本??车（不是什么爱过情怀）心里作用 别喷！最后叫朋友到处看车 1.第一次看的是长安逸动 价格是便宜 基本上有的功能还是有 无赖没有esp气囊有点少 外形还不错 暂定。2.起亚k4和新k3 k4还不错 就是价格超出预算 也没用购置税减半！pass了 k3就我感觉就很一般了。3.比亚迪思锐:车是好车 配置也挺不错 可惜已经停产 4 比亚迪宋:外观配置真没的说 考虑到2.0t油耗大 以后维修成本高 城市道路还是自吸的好 预算也超了 5 吉利新帝豪 外观配置还行！暂定！6 陆风x5plus|改款新车 国产配置真没的说 老款x5看论坛口碑真不怎么好 生锈 芭蕉熟了之类的 只能先pass了！其他就不细细说了 看了挺多的 科鲁兹 c4 408等等！后来买领动是我最开始看到小区里好多elantra这车 百度下是伊兰特 最后看帖子才知道是朗动 加上快上市的领动就是4代同堂了！上之家看了下价格预算内 叫上朋友直接去4s店看朗动 各方面都不错 也挺好看的 除了车头有点短外 口碑也还不错！最后都准备订了！可以看我前面的帖子！最后看到领动外形比朗动还好看 问了几个销售都说在名图和朗动之间 估计12w起！价格还不确定 我更喜欢领动 考虑到买车不用着急 等等领动上市！上市第2天就出配置了 看了基本上够用 也有esp 第3天就跑到4儿子店去问了！去的太早还不知道有没有免息活动也不知道能不能加选装3 就和4s约定如果不能加装3和没有免息活动就改朗动自尊！选装3装逼点 谈好送的 交定金 走人等消息！4月1号那天接到4s电话说可以加装3 没有免息 考虑到更喜欢领动 再者新车更新换代 和老婆商量了下打算全款！给4s去电话就算选定领动了 坐等提车！14号那天接到电话说车到了 家里人觉得购车也是这么大一笔开支 得看个日子去提 选定19号（农历3月13 初3 13 23太上老君3不管 意思代表日子不错） 没办法老人家的想法也得尊重下！！！！！！前面话太多了 价格和送的东西我后面再细说 各位看官见谅 说了这么多直接上图！4儿子店展车提车看了下发动机有无其他异响 我就是小白一个 叫朋友听听声音的提车时的公里数检查完毕 交钱 上保险 打临牌上路加油咯！第一顿得吃饱点才有劲 也可以看看有没有漏油 也可以听听开车时油箱有没有撞击声远看 还是挺不错的正前 大气不自带导航 不过有carplay和carlife连手机 地图更新更快哦！中控还是挺好看的 个人比较喜欢?? 自己喜欢几天 何必在意别人的想法呢！  [1] [2] [3] [4] [5] [下一页]"|http://www.qc188.com/czsc/201605/131821.html|2016-05-23
기타|2457720372|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-23 14:17:06|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=126&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-23
其他媒体|2457767157|zhidao_baidu|东芝|ZHO|2016-05-23 14:44:02|东风悦达起亚k3高配全款多少钱曲阳4s店|汽车东风悦达起亚k3高配全款少钱曲阳4s店|http://zhidao.baidu.com/question/2055587863683453427.html?fr=qlquick&entry=qb_list_default|2016-05-23
기타|2457816663|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 15:12:05|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=107&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2457816896|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 15:12:06|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=63&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-23
기타|2457831966|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-23 15:23:16|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=219&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-23
기타|2457863901|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 15:40:04|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=118&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2457864193|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 15:40:05|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=47&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-23
기타|2457877245|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 15:46:04|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=108&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2457877373|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 15:46:04|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=64&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-23
기타|2457879407|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-23 15:47:14|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=130&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-23
기타|2457890856|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-23 15:54:02|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=222&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-23
기타|2457891244|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-23 15:54:03|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=69&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2457925855|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 16:12:02|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=48&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-23
기타|2457934791|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-23 16:17:48|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=132&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-23
기타|2457992942|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 16:47:29|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=120&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2457993073|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 16:47:29|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=50&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-23
기타|2457993841|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 16:47:30|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=109&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2457993890|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 16:47:30|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=65&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-23
기타|2458003579|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-23 16:52:02|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=134&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-23
기타|2458019324|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-23 17:00:06|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=71&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2458052470|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 17:20:07|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=121&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2458066236|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-23 17:25:02|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=135&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-23
기타|2458100905|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-23 17:43:01|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=114&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-23
기타|2458105949|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 17:45:04|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=51&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-23
기타|2458121001|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 17:52:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=110&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2458121178|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 17:52:01|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=66&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-23
기타|2458211073|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 18:41:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=123&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2458211242|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 18:41:01|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=53&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-23
기타|2458235228|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 18:54:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=111&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2458235376|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 18:54:01|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=67&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-23
기타|2458259806|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-23 19:07:29|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=115&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-23
기타|2458312123|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-23 19:39:02|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=116&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-23
기타|2458329378|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 19:49:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=124&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2458329565|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 19:49:03|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=54&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-23
기타|2458331559|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 19:50:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=113&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2458331709|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 19:50:03|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=69&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-23
기타|2458336059|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-23 19:53:01|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=136&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-23
기타|2458417238|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-23 20:43:01|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=117&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-23
기타|2458446098|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-23 20:58:02|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=223&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-23
기타|2458449299|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-23 21:00:01|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=138&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-23
기타|2458494137|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 21:27:43|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=71&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-23
기타|2458494606|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-23 21:27:50|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=141&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-23
기타|2458499561|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-23 21:30:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=225&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-23
기타|2458552250|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-23 22:01:03|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=74&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2458560876|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 22:06:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=115&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2458608772|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-23 22:35:02|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=142&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-23
기타|2458651285|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 22:59:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=125&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2458660778|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-23 23:05:01|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=144&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-23
기타|2458683590|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 23:20:14|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=116&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2458684938|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-23 23:21:03|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=72&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-23
기타|2458705717|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-23 23:30:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=75&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2458710672|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 23:33:12|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=127&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-23
기타|2458711671|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-23 23:34:01|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=57&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-23
기타|2470070169|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 00:05:01|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=81&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-30
기타|2470103317|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 00:34:05|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=209&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2470103408|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 00:34:05|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=140&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-30
기타|2470444898|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 08:04:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=210&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2470474935|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 08:38:03|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=141&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-30
기타|2470476907|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 08:39:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=82&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-30
기타|2470562357|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 09:51:01|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=100&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-05-30
기타|2470562402|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 09:51:01|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的。....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=82&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-05-30
기타|2470562408|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 09:51:01|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=79&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-05-30
各大媒体|2470793025|12365auto|质量投诉|ZHO|2016-05-30 12:07:20|东风悦达起亚K3经销商欺骗客户卖库存车|投诉编号：【142205】 投诉品牌： 东风悦达起亚 投诉车系： 起亚K3 投诉车型： 2015款 1.6L 手动 GLS 投诉时间： 2016-05-28 17:43    投诉内容： 我在2015年11月29日早上大约十点去的店 在中午两点左右选好车 三点左右谈好价格 在后面的过程中 我给他们说我要现车 还要求不要库存车 他们给我回答的是他们店没有库存车 都不超过三个月 然后我说我全款今晚要提车 再后面他们让我等 大概四点半左右 他们开出来一辆白的k3我说车是什么时候他们说2015年7月份的 我说超了3个月 他们就给我解释说从江苏运过来要两个月 在他们这儿放了2个月左右 我害怕他们弄错问了好多次 因为他们快下班了 他们开始让我交钱 我的车价是102000我付清了 但发票他们打了98000接着他们催促我给他们的服务态度做个评价 我就签了名 在交钱是钱了个名 合同自始至终没见到 我弄完五点半了 他们要下班 说手续邮给我 我就开车回家了 直到一月份我挂完牌子 我朋友发现我的车2014年7月份的 我立马回家给销售顾问打电话 他还在骗我说我的车是2015年7月的 不不算车门 要看合格证上的 并且给我承诺是2014年7月份的话要满足我提的要求 这个通话有录音 我回家看了合格证也是2014年7月的 我联系销售顾问 他说我自认倒霉把 给厂家打电话 他们先是说给我处理 一个月以前又说他们也没办法 唉 我是个老师 钱存了买个车 就成了这样 为什么我们这些人去哪里都被欺负 像这些4s店 人随便骗 发票可以乱打 真的是无法无天吗？为什么咱们国家的市场这么乱 社会氛气这么差 唉。   投诉回复： 车质网已将您的投诉转给生产企业以及政府有关主管部门 我们将会对此投诉继续跟踪 请您持续关注！|http://www.12365auto.com/zlts/20160528/142205.shtml|2016-05-30
기타|2470834920|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 12:36:14|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=179&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2470835363|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 12:36:14|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=135&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-30
기타|2470880997|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-30 13:01:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=121&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2470889900|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 13:06:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=181&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2470889951|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 13:06:02|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=137&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-30
기타|2470943057|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 13:40:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=180&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2470943124|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 13:40:02|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=136&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-30
기타|2471032891|Autohome_review|랑동(朗动)|ZHO|2016-05-30 14:35:01|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=187&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-30
기타|2471045762|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 14:42:02|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=183&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-05-30
기타|2471046016|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 14:42:03|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=101&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-05-30
기타|2471046081|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 14:42:03|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的。....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=83&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-05-30
기타|2471046089|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 14:42:03|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=80&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-05-30
기타|2471061483|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-30 14:51:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=122&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471069385|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-30 14:55:02|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=157&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-30
기타|2471102629|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 15:15:05|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=182&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471103329|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 15:16:08|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=138&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-30
其他媒体|2471137041|zhidao_baidu|电子数码 > 手机/通讯-手机使用|ZHO|2016-05-30 15:34:01|本田凌派 起亚k3'标志308'大众朗逸 丰田雷凌！谁更值得拥有 请说明理由 由于本人对车不太了解|汽车丰田由于本人对车不太了解;标志308' 起亚k3' 买个车也不容易 我不想让自己太后悔 丰田雷凌;大众朗逸 请说明理由！谁更值得拥有本田凌派|http://zhidao.baidu.com/question/1434260605162465019.html?fr=qlquick&entry=qb_list_default|2016-05-30
기타|2471140348|Autohome_review|랑동(朗动)|ZHO|2016-05-30 15:36:02|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=191&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-30
기타|2471145155|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 15:38:14|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=211&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471145348|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 15:38:15|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=142&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-30
기타|2471145522|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 15:38:15|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=83&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-30
기타|2471152617|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 15:43:02|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=186&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-05-30
기타|2471152888|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 15:43:09|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=104&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-05-30
기타|2471152934|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 15:43:10|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的。....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=86&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-05-30
기타|2471152944|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 15:43:10|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=83&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-05-30
기타|2471164436|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-30 15:49:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=127&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471248150|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 16:36:06|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=215&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471248424|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 16:36:06|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=146&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-30
기타|2471248818|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 16:37:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=86&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-30
기타|2471262491|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 16:43:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=184&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471262544|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 16:43:02|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=140&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-30
기타|2471286232|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-30 16:55:02|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=158&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-30
기타|2471305899|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 17:07:30|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=216&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471306163|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 17:07:30|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=147&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-30
기타|2471306428|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 17:07:35|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=87&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-30
기타|2471321014|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 17:17:32|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=185&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471321384|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 17:18:14|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=141&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-30
기타|2471349259|Autohome_review|랑동(朗动)|ZHO|2016-05-30 17:30:02|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=192&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-30
기타|2471360474|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 17:37:01|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=187&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-05-30
기타|2471362505|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 17:38:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=88&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-30
기타|2471393482|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-30 17:53:03|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=128&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471464965|Autohome_review|랑동(朗动)|ZHO|2016-05-30 18:31:01|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=194&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-30
기타|2471474251|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 18:36:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=219&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471474465|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 18:36:06|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=150&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-30
기타|2471474601|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 18:36:06|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=90&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-30
기타|2471479544|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 18:39:02|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=189&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-05-30
기타|2471479781|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 18:39:02|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=107&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-05-30
기타|2471479830|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 18:39:02|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的。....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=89&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-05-30
기타|2471479837|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 18:39:02|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=86&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-05-30
기타|2471516573|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 18:59:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=187&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471516739|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 18:59:02|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=143&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-30
기타|2471563693|Autohome_review|랑동(朗动)|ZHO|2016-05-30 19:27:52|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=196&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-30
기타|2471575192|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 19:34:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=218&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471575317|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 19:34:01|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=149&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-30
기타|2471599637|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-30 19:49:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=129&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471667987|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 20:30:04|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=91&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-30
기타|2471694534|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-30 20:45:03|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=130&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471696638|Autohome_review|랑동(朗动)|ZHO|2016-05-30 20:46:01|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=197&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-30
기타|2471769339|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 21:31:02|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=190&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-05-30
기타|2471769564|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 21:31:02|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=108&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-05-30
기타|2471769591|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 21:31:02|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的。....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=90&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-05-30
기타|2471769594|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 21:31:02|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=87&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-05-30
기타|2471794762|Autohome_review|랑동(朗动)|ZHO|2016-05-30 21:46:02|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=198&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-30
기타|2471806621|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 21:53:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=191&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471806736|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 21:53:02|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=146&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-30
기타|2471860010|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 22:27:34|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=221&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471860105|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 22:27:34|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=152&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-30
기타|2471882162|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-30 22:40:03|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=133&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471902377|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 22:52:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=192&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471902472|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 22:52:02|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=148&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-30
기타|2471908063|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 22:56:01|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=93&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-30
기타|2471951991|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 23:24:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=193&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471952140|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-30 23:24:01|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=149&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-30
기타|2471957758|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 23:27:48|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=222&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-30
기타|2471957876|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 23:27:48|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=153&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-30
기타|2471961129|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 23:29:01|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=191&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-05-30
기타|2471961348|Autohome_review|K3(起亚K3)|ZHO|2016-05-30 23:29:02|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=109&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-05-30
기타|2472003294|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-30 23:56:04|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=94&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-30
기타|2504028076|Autohome_review|K3(起亚K3)|ZHO|2016-06-17 01:08:01|2016年06月16日 发表了口碑|来自：汽车之家Android版  2016年06月16日 发表了口碑  口碑   《用车差不多一个月 对K3还是挺满意挺喜欢的。》           【最满意的一点】第一是外形 实车比相片好看多了。【最不满意的一点】扶手箱比较短 又不能前后移动。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】因为我是个韩国迷 很多韩剧都是用起亚车代言 所以很喜欢 这车我自己也试驾过很多次（因为有亲戚在起亚4S店工作 k3的行车隔音比凌派好 动力又比福睿斯 轩逸 等等要强。买K3之前我考虑过雷凌 朗逸 雷凌的外形我挺喜欢的 CVT无级变速器的行驶平顺性曾经让我很喜欢 但是比K3贵 所以不要 朗逸确实是很不错 开起来很舒服 底盘对于一些小颠簸过滤的很好 朗逸真的挺好 不过还是比K3贵 空间也没有K3大。【其他描述】|http://k.autohome.com.cn/spec/19724/view_1167733_1.html?st=8&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2504119115|Autohome_review|K3(起亚K3)|ZHO|2016-06-17 02:23:03|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=196&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2504119149|Autohome_review|K3(起亚K3)|ZHO|2016-06-17 02:23:03|2016年05月19日 发表了质量评价|2016年05月19日 发表了质量评价  质量   【行驶过程】  刹车时有异响-车辆前部  【内饰】  随车脚垫会滑动或污损       来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=179&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2504119153|Autohome_review|K3(起亚K3)|ZHO|2016-06-17 02:23:03|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=176&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2504119295|Autohome_review|K3(起亚K3)|ZHO|2016-06-17 02:23:03|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=88&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2504119326|Autohome_review|K3(起亚K3)|ZHO|2016-06-17 02:23:03|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=74&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2504119366|Autohome_review|K3(起亚K3)|ZHO|2016-06-17 02:23:03|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=52&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2504119502|Autohome_review|K3(起亚K3)|ZHO|2016-06-17 02:24:01|2016年06月16日 发表了口碑|来自：汽车之家Android版  2016年06月16日 发表了口碑  口碑   《用车差不多一个月 对K3还是挺满意挺喜欢的。》           【最满意的一点】第一是外形 实车比相片好看多了。【最不满意的一点】扶手箱比较短 又不能前后移动。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】因为我是个韩国迷 很多韩剧都是用起亚车代言 所以很喜欢 这车我自己也试驾过很多次（因为有亲戚在起亚4S店工作 k3的行车隔音比凌派好 动力又比福睿斯 轩逸 等等要强。买K3之前我考虑过雷凌 朗逸 雷凌的外形我挺喜欢的 CVT无级变速器的行驶平顺性曾经让我很喜欢 但是比K3贵 所以不要 朗逸确实是很不错 开起来很舒服 底盘对于一些小颠簸过滤的很好 朗逸真的挺好 不过还是比K3贵 空间也没有K3大。【其他描述】|http://k.autohome.com.cn/spec/19724/view_1167733_1.html?st=9&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-17
其他媒体|2504488639|zhidao_baidu|文化/艺术|ZHO|2016-06-17 09:41:04|东风悦达起亚k3摇控器放在车里怎样打开车门|汽车|http://zhidao.baidu.com/question/266441291454531845.html?fr=qlquick&entry=qb_list_default|2016-06-17
기타|2504784694|Autohome_review|K3(起亚K3)|ZHO|2016-06-17 12:45:03|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=193&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2504784729|Autohome_review|K3(起亚K3)|ZHO|2016-06-17 12:45:03|2016年05月19日 发表了质量评价|2016年05月19日 发表了质量评价  质量   【行驶过程】  刹车时有异响-车辆前部  【内饰】  随车脚垫会滑动或污损       来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。还有它的外形吧 .【最不满意的一点】买的自动挡的 动力比较弱 起步和超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 在高速上声音很大.隔音也不咋地啊. 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】虽然比较喜欢老款.虎啸脸.新款改了前脸进气格栅 但看着也是挺大气的.韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 宝俊560亲戚家有一辆了 不想买一样的 哈弗H6确实好看 就怕发动机不给力啊 本来就打算定福睿斯了 期间也看了好多次了 51和姐夫一起去车展看福睿斯的 销售特别的热情 姐夫比较懂车 看了看说福睿斯 觉得不咋地 说屁股太丑 要不然在考虑考虑 然后又转了几圈 走到了起亚的展台 看到了16款的k3还不错 我以前只是偶尔关注过起亚 对它了解不是很多 正好我姐夫的朋友前几天买了一台k3.优惠还行.我就问了一下还有没有老款的 销售说老款的卖完了只有新款的了 但是我还是觉得老款的看着大气 新款看着比较秀气 仔细想想这个价位的车都差不多 主要功能就是家庭代步 就和销售砍价 因为是51车展 所以优惠比较大 本来想分期买的 因为没有房贷什么的 压力不是很大 而且分期还能多送个导航 但是分期需要的手续太麻烦 老爸说那就全款吧 然后就定了k3 事后我在之家上面了解到销售给我的优惠还是挺大的啊 比心理预期的好点.因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的啊。.....|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=176&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2504784742|Autohome_review|K3(起亚K3)|ZHO|2016-06-17 12:45:04|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=173&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2504784876|Autohome_review|K3(起亚K3)|ZHO|2016-06-17 12:45:04|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=85&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2504784896|Autohome_review|K3(起亚K3)|ZHO|2016-06-17 12:45:04|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=71&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2504784921|Autohome_review|K3(起亚K3)|ZHO|2016-06-17 12:45:04|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=49&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2504805982|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-17 13:00:01|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=69&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2504892161|Autohome_review|BYD S6(比亚迪S6)|ZHO|2016-06-17 13:59:01|2016年04月01日 发表了口碑|来自：汽车之家iPhone版  2016年04月01日 发表了口碑  口碑    《空间大就不用说了 没有之前担心的动力不足 感觉动力够用》           【最满意的一点】空间 配置 虽然2.0手豪（不想要天窗 应人而异）但是后期选装自装也是感觉很霸气 好多十多万的车都没有的配置  心里美滋滋～【最不满意的一点】目前就发现右后轮起步有点异响 但是说来也怪  每次到4s店就没有了 去了四五次都不响了 回家没几天又继续  好邪～【空间】前几天去了东北  （有贴） 后面气垫床谁俩人（178cm）没问题  还能装点东西～【动力】没有网上说的那么肉  我只想说只要舍得给油什么车都不肉【操控】开的还不错  就是刚开始开离合太高不习惯  现在习惯了 感觉很透  油门也挺灵活  （之前在部队开猛士） 开小六感觉 很棒【油耗】比预计要低可能跑长途的 以前市区差不多9个油还能接受 这次高速回来平均降到8.7 不管多少2.0这么大的车 只要不超十个油都能接受【舒适性】椅子倍舒服 以前猛士没法比  也不能比 不是一个级别 感觉比朋友的k3舒服多了！【外观】外观挺不错的  不过现在出来好的新车自然小六要逊色不少  不过自己折腾加装踏板 牛头杠 行李架 （准备换Q5大灯和仿宝马LED尾灯）【内饰】内饰除了座椅和方向盘很满意 其他都很一般般吧！【性价比】性价比就不说了直接满分  这么大的车裸车7w多块钱 去哪找？【为什么最终选择这款车？】其实购车前一直看中h6  但是资金有限（不想贷款）全身就10w  后来看了好多款  家里差点让买了宝骏560  和陆丰x7（家里支持资金）但是最后还是选择了s6 因为家里不喜欢比亚迪 这个名字（大家好多都懂的）说十几万宁愿买个CRV  不过我不喜欢日产（还是应人而异）【其他描述】|http://k.autohome.com.cn/spec/18563/view_1041472_1.html?st=193&piap=0 2088 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2504899787|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-17 14:03:07|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=70&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2505020894|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-17 15:21:21|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=72&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-17
其他媒体|2505041804|zhidao_baidu|电脑/网络 > 硬件 > 显示器|ZHO|2016-06-17 15:34:01|东风悦达起亚k3漳浦哪一家卖|汽车汽车购买东风悦达起亚k3漳浦哪一家卖|http://zhidao.baidu.com/question/1641774840014612500.html?fr=qlquick&entry=qb_list_default|2016-06-17
기타|2505108075|315che|行情|ZHO|2016-06-17 16:14:43|2016款起亚K3降价促销 现金直降售全国|　　【天津行情】近日 中国汽车消费网编辑走访获悉 北京仁祥宏业4s店内起亚K3现车销售 颜色可选 目前购车部分车型可优惠5万元 感兴趣的朋友可以到店咨询购买 厂家的活动价格促销 当天可提走现车 没有任何附加条件 希望诚心购买人士到店详谈。详情请拨起亚/K3销售热线:*********** 刘经理 以下是2015款起亚K3的具体的报价表：北京地区起亚最新价格：起亚K3报价表（2016-06-17）车型指导价销售价优惠情况现车情况起亚K3 2015款 1.6L MT GL10.28万5.28万5万现车充足起亚K3 2015款 1.6L AT GL11.28万6.28万起亚K3 2015款 1.6L AT GLS12.48万7.48万起亚K3 2015款 1.6L AT DLX13.18万8.18万起亚K3 2015款 1.6L AT Premium14.38万9.38万起亚K3 2015款 1.8L AT Premium14.98万9.98万中国汽车消费网制表　　起亚K3各地行情信息请关注：http://auto.315che.com/qiyak3/articles__43.htm　　更多同级别车型价格变动信息请关注：http://www.315che.com/hq/　　基本介绍：2015款K3的前中网颜色变更 后保险杠和排气管也经过了重新设计 DLX AT及以上车型配备了椭圆形的镀铬排气管。2015款K3还新增珍珠白这一可选车身颜色。中控面板位置的空调按钮增加镀铬装饰 车内引入了更多软性材料装饰。2015款K3的主要竞争对手还是目前市场上主流的紧凑型轿车 例如现代朗动、本田凌派、雪佛兰科鲁兹等。和竞争对手相比 丰富的配置和个性的造型是吸引不少消费者选择K3的因素。  起亚K3 指导价： 10.28～14.98 万   品牌：起亚图片(共767 张)   配置   车吧   报价   口碑(共133 条)315che.com 　　配置详解：GL配备了主副驾驶座安全气囊、ABS+EBD、多功能方向盘上下调节、行车电脑显示屏、前座中央扶手、前雾灯、大灯高度可调、后视镜电动调节、后视镜加热、手动空调。　　GLS多了日间行车灯、后排杯架、后座中央扶手、座椅高低调节、真皮方向盘、电动天窗、无钥匙启动系统以及选装配置倒车视频影像、真皮座椅、腰部支撑调节、前排座椅电动调节、电动座椅记忆、座椅通风、GPS导航系统、蓝牙/车载电话等。　　DLX在GLS的基础上又多了EBD+EBA+ASR、真皮座椅、后座出风口和温度分区控制。　　Premium作为最高配 新增了后视镜电动折叠、后视镜记忆、氙气大灯、电动座椅记忆、前排座椅加热、座椅通风、前排座椅电动调节、腰部支撑调节、方向盘换挡、定速巡航、胎压监测装置。自动挡还可选装前/后排头部气囊(气帘)。　　注：中国汽车消费网 (www.315che.com) 提供的价格信息为编辑采集的及时信息 价格仅供参考 车市行情天天变 消费者如需购买相关车型 应该尽快与具体经销商电联或当面洽谈。另 文中引用图片和推荐经销商仅为资料信息 与价格信息来源无关。|http://inf.315che.com/n/2016_06/689439/|2016-06-17
기타|2505143203|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-17 16:33:01|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=74&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2505191368|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-17 17:00:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=215&piap=0 78 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2505267539|Autohome_review|아반떼 AD(领动)|ZHO|2016-06-17 17:44:03|2016年06月02日 发表了口碑|来自：手机汽车之家  2016年06月02日 发表了口碑  口碑    《外观拉风 配置足够 整体性价比还是不错的。》           【最满意的一点】外观很拉风 现在路上还很少见 大轮毂。日间行车灯很高大上 自动头灯也很高端。中控台是软的 车内显示屏清晰度很高。倒车影像有随动辅助导线。很方便。车内音响很赞 我喜欢听音乐 完全满足我的要求。【最不满意的一点】后排不能放倒 这个真心很郁闷 这个放倒真的很难吗？这几天B柱内有异响 这还是新车呀 哎。。过几天去4s看看 希望不是啥大问题。另外胎噪确实大 我想跟轮胎大也有关系吧。悬挂还是有点硬 不过在接受范围内。【空间】空间同级别还是有优势的 中间无凸起。【动力】动力够用 现在用的eco模式【操控】转向精准 没啥虚位。【油耗】表显6 肯定是不准的 等下次油表亮再算算。【舒适性】还可以 家用够了。【外观】满意【内饰】做工还是比较好的 接缝均匀。【性价比】性价比高【为什么最终选择这款车？】同级别都看了 也试驾了 福克斯空间太小 科鲁兹都说油耗高 新英朗有点老气 卡罗拉没esp 思域根本没现车 看来看去家用也就韩系车了。【其他描述】换车的想法去年就有了 但是一直没有付诸行动 一是因为暂时有车开 二是今年上市新车多 想再等等 经常看论坛 心里已经有了几个备选 英朗 老表刚买的 开始觉得性价比很高 后来发现新旧差别很大 就pass了。福克斯外观不错 但是同事有好几辆 不想买一样的。k3性价比很高 优惠很大 但是新款感觉你没老款好看。看到最后就是领动了 配置高 外观拉风 总体性价比很高。|http://k.autohome.com.cn/spec/25701/view_1148059_1.html?st=52&piap=0 3959 0 0 2 0 0 0 0 0 1|2016-06-17
其他媒体|2505282973|bitauto|易车 > 问答 > 问题分类|ZHO|2016-06-17 17:53:01|东风悦达起亚k31·；4t发动机|东风悦达起亚k31·；4t发动机     提问者：易车网友 分类：  东风  买车  汽车知识  浏览[4]  2016-06-17 16:46  举报   东风悦达起亚k31·4t发动机|http://ask.bitauto.com/detail/6673639/?leads_source=p029001|2016-06-17
기타|2505293334|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-17 18:00:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=216&piap=0 78 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2505370015|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-06-17 18:46:04|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=217&piap=0 78 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2505426641|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-17 19:19:02|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=77&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2505465603|Autohome_review|잉랑GT(英朗)|ZHO|2016-06-17 19:45:02|2016年06月12日 发表了口碑|来自：手机汽车之家  2016年06月12日 发表了口碑  口碑   《颜值尚佳 空间大方 配置丰富 油耗满意 性价比高。》             【最满意的一点】外形没得说大家都说好看 空间大老妈坐了说不会头晕很舒服 静音效果还行。【最不满意的一点】冷车启动发动机有点抖动 喇叭滴滴声小气 悬挂有点硬 加速不够平顺 漆面有点薄 动力凑合用。【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】看的可多了都有丰田卡罗拉（没ESP）起亚k3（换前脸了）现代朗动（领动上市）现代领动（优惠少）马自达昂科赛拉（后排空间太小了）别克新英朗（标配ESP 直瀑前脸 侧线条刚毅 油耗适中 空间很大 优惠不错）懂你说的 懂你没说的 各项指标均匀 值得拥有。【其他描述】|http://k.autohome.com.cn/spec/25864/view_1159235_1.html?st=78&piap=0 982 0 0 2 0 0 0 0 0 1|2016-06-17
기타|2521793127|Autohome_review|랑동(朗动)|ZHO|2016-06-27 00:00:01|2016年06月21日 发表了口碑|来自：手机汽车之家  2016年06月21日 发表了口碑  口碑   《外观时尚好看 车子配置高实惠》           【最满意的一点】车子的外观和空间【最不满意的一点】1.6发动机动力不足【空间】后排虽然不能放倒 但足够日常生活所用 如何是放大东西的话就放不进去了【动力】起步肉 加速平稳 如果跑高速的话 油门响应有点慢 比如在跑高速过程中 你松下油门再想加速踩油门要踩深一点 中间有2秒的停顿加速【操控】方向盘轻 方向比较准【油耗】综合油耗还可以接受【舒适性】座椅很舒服 胎噪比较大跑高速【外观】外观非常喜欢【内饰】内饰中控台是软的比思域硬胶好很多【性价比】配置高 价格便宜实惠【为什么最终选择这款车？】选车中看了思域 速腾 卡罗拉 雷凌 k3。朗动的外观内饰价格优惠吸引我【其他描述】|http://k.autohome.com.cn/spec/20618/view_1178572_1.html?st=30&piap=0 2764 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2521916980|Autohome_review|닛산 티아나(天籁)|ZHO|2016-06-27 01:35:03|2016年06月20日 发表了口碑|来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《性价比超高 外观大气稳重 省油。》             【最满意的一点】坐椅舒适 减震不错 空间宽敞 电动坐椅 后排出风口非常好。【最不满意的一点】自动大反应慢 基本没用 舒适版无倒车雷达 好歹十几万的车 居然不配这个两百块钱又非常实用的东西？前保险杠与叶子板接合处是水平状态 下雨天开车后污垢会从接合处流到保险杠上 很难看 我观察过其他车 其他车的这个部位一般都是有一个角度的 污水会顺着角度流到地上 不会弄脏保险杠 我认为这是设计不到位。【空间】很满意 现在看别人家的车都觉得小【动力】比原来的1.4强多了。【操控】没开过其他车 反正比k2好【油耗】没k2省 不过排量大0.6车重四百公斤 很不错了。我最低开过3.6升百公里 一般来说两百块跑四百三四十公里 高速城区农村各有一部分 如果纯城区只能跑三百六十左右。【舒适性】不错 买天籁就是冲这个来的 我腰椎间盘突出 做了手术 上了钢筋的 不能受冲击 过减速带比原来好多了【外观】大气稳重【内饰】还行 有味 但比原车好。【性价比】超高 别人都说这车得二十几万吧 我说十五万没人信。【为什么最终选择这款车？】由于前一个车是起亚k2 所以最先看的是k3 媳妇试坐之后认为除了大点之外和k2没啥区别 后来又试了一些其他车 都没感觉 直到走进一家店里看到天籁 媳妇坐进去试了一下 感觉很满意 移沙发确实不错 但是就是觉得价格超了 那是去年的事了 今年三月又去试了kx3 板车悬挂同样让人不满意 本地车展又去转了转 带媳妇去看了丰田卡罗拉 内饰丑死个人 比老款难看多了 后来媳妇发话 干脆一步到位 上天籁。【其他描述】|http://k.autohome.com.cn/spec/15104/view_1173431_1.html?st=47&piap=0 634 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2521935844|Autohome_review|포커스(福克斯)|ZHO|2016-06-27 01:51:02|2016年06月20日 发表了口碑|"来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《唯一缺点就是空间小！》           【最满意的一点】好开 很稳 很省心 【最不满意的一点】空间小 降价快【空间】坐五个人不是太挤 后备箱比较大 综合还是不错【动力】不开空调 一个人开还是不错的 要舍得给油！驾驶乐趣不错 满座来空调那就力不从心了【操控】转向精准 悬架支撑不错 过弯比较有信心 过坑洼路面不是太舒服！【油耗】油耗还能接受 不是太高！当然没发和日系车比咯！【舒适性】座椅包裹性好 不过长途驾驶感觉不太舒服 座椅不是太软。关窗静音效果不错 胎噪有点大 其他方面都还不错的！【外观】外观还是比较漂亮的！轮毂再大一号就帅多了！【内饰】用料不错 做工就不敢恭维了！缝隙太大 不像合资的车。哎！真是应征了网友们所说的?百年福特毁于长安！希望长安福特之后们在做工方面改善改善！【性价比】性能不错 安全配置比较齐全 长安的价格贬值比较快！很让消费者伤心??买了车快两年了 唯一后悔的就是不该买最低配版的 如果再给我重新选择的机会 毫不犹豫直接上中高配！！！！！！！！！！【为什么最终选择这款车？】朗动 k3|朗逸。朗动挺漂亮 老婆看的时候说感觉太单薄.k3和朗动差不懂 配置也差不多 朋友的也是k3|不想大家都买一样的 果断放弃。朗逸神车 比较中庸 保值率高 不适合我们九零后 要有个性。福克斯基本安全配置比较高 油耗必上一代有所改善 车身扎实。比较适合自己 空间勉强够用 主要是自己开 能接受。【其他描述】油箱负压 空调效果不是很好 保养贵"|http://k.autohome.com.cn/spec/12132/view_1176643_1.html?st=103&piap=0 364 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522097957|Autohome_review|랑동(朗动)|ZHO|2016-06-27 05:53:02|2016年06月21日 发表了口碑|来自：手机汽车之家  2016年06月21日 发表了口碑  口碑   《外观时尚好看 车子配置高实惠》           【最满意的一点】车子的外观和空间【最不满意的一点】1.6发动机动力不足【空间】后排虽然不能放倒 但足够日常生活所用 如何是放大东西的话就放不进去了【动力】起步肉 加速平稳 如果跑高速的话 油门响应有点慢 比如在跑高速过程中 你松下油门再想加速踩油门要踩深一点 中间有2秒的停顿加速【操控】方向盘轻 方向比较准【油耗】综合油耗还可以接受【舒适性】座椅很舒服 胎噪比较大跑高速【外观】外观非常喜欢【内饰】内饰中控台是软的比思域硬胶好很多【性价比】配置高 价格便宜实惠【为什么最终选择这款车？】选车中看了思域 速腾 卡罗拉 雷凌 k3。朗动的外观内饰价格优惠吸引我【其他描述】|http://k.autohome.com.cn/spec/20618/view_1178572_1.html?st=32&piap=0 2764 0 0 2 0 0 0 0 0 1|2016-06-27
其他媒体|2522216275|zhidao_baidu|电子数码 > MP4/MP3|ZHO|2016-06-27 08:43:02|东风悦达起亚k3码数拉不上怎么回事|汽车东风悦达起亚k3码数拉不上怎么回事|http://zhidao.baidu.com/question/2205675317323665068.html?fr=qlquick&entry=qb_list_default|2016-06-27
기타|2522253252|Autohome_review|닛산 티아나(天籁)|ZHO|2016-06-27 09:17:01|2016年06月20日 发表了口碑|来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《性价比超高 外观大气稳重 省油。》             【最满意的一点】坐椅舒适 减震不错 空间宽敞 电动坐椅 后排出风口非常好。【最不满意的一点】自动大反应慢 基本没用 舒适版无倒车雷达 好歹十几万的车 居然不配这个两百块钱又非常实用的东西？前保险杠与叶子板接合处是水平状态 下雨天开车后污垢会从接合处流到保险杠上 很难看 我观察过其他车 其他车的这个部位一般都是有一个角度的 污水会顺着角度流到地上 不会弄脏保险杠 我认为这是设计不到位。【空间】很满意 现在看别人家的车都觉得小【动力】比原来的1.4强多了。【操控】没开过其他车 反正比k2好【油耗】没k2省 不过排量大0.6车重四百公斤 很不错了。我最低开过3.6升百公里 一般来说两百块跑四百三四十公里 高速城区农村各有一部分 如果纯城区只能跑三百六十左右。【舒适性】不错 买天籁就是冲这个来的 我腰椎间盘突出 做了手术 上了钢筋的 不能受冲击 过减速带比原来好多了【外观】大气稳重【内饰】还行 有味 但比原车好。【性价比】超高 别人都说这车得二十几万吧 我说十五万没人信。【为什么最终选择这款车？】由于前一个车是起亚k2 所以最先看的是k3 媳妇试坐之后认为除了大点之外和k2没啥区别 后来又试了一些其他车 都没感觉 直到走进一家店里看到天籁 媳妇坐进去试了一下 感觉很满意 移沙发确实不错 但是就是觉得价格超了 那是去年的事了 今年三月又去试了kx3 板车悬挂同样让人不满意 本地车展又去转了转 带媳妇去看了丰田卡罗拉 内饰丑死个人 比老款难看多了 后来媳妇发话 干脆一步到位 上天籁。【其他描述】|http://k.autohome.com.cn/spec/15104/view_1173431_1.html?st=48&piap=0 634 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522345228|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 10:23:11|2016年06月18日 发表了口碑|"2016年06月18日 发表了口碑  口碑    《空间大 省油 外观大气 优惠力度大》             【最满意的一点】空间大 油耗低 外观时尚 1万公里换机油保养。【最不满意的一点】没有ESP 没有发动机防盗 这俩项确实不应该简配。【空间】买车前参考过昂克赛拉 起亚k3|朗动 轩逸 蓝鸟 朗逸。轴距都是2700mm|但是看罗拉空间明显要大一些。180的大长腿坐进去都不挤。后排地面中间平整 也没有扶手 座三个175的壮汉也不觉得挤 不过后备箱不如轩逸的 感觉略小。【动力】1.6L的动力一个人开经常会有推背感 毕竟122马力 哈哈 但是座人了就感觉肉了 不过比朋友的斯柯达明锐1.6L双离合还是强劲不少 而且自然吸气的发动机跟涡轮增压比起来也没有烧机油的风险。【操控】之前开过面包车 开过荣威 但是跟卡罗拉的CVT比起来差远了 卡罗拉的标定确实比较扎实 换挡逻辑非常清新 开起来很平顺 出乎意料。在市区基本在1000转左右 处于ECO模式 高速跑120迈也就不到2000转左右 不知道需不需要像有的老司机说的过了磨合期高速拉缸。【油耗】刚提车时候油耗归零 开了110公里 竟然达到了惊人的4.1L/百公里 后来随着里程的增加逐步稳定在了6.5 6.6。日系车省油的名号确实不是盖的。【舒适性】这个价位的卡罗拉没有独立悬挂确实有些遗憾 在过减速带的时候 感觉略硬 风噪没有群友说的夸张 到了100迈内部还是比较安静的 但是偶尔能听到像石子刮地的声音 一直找不到原因。【外观】外观比老款的确实好看 个人觉得比雷凌的要收敛 离地间隙很低 好看但是也容易被磕碰。【内饰】内饰是硬塑料 黑白小仪表。10寸导航很加分 很大气 堪比K3.织物座椅去淘宝配个坐垫 美观舒适 朋友的真皮座椅夏天烫屁股。置物空间很多 放置杂物什么的没问题。【性价比】恰逢五一车展搞活动 优惠力度还是比较大了 送了贴膜导航装具行车记录仪。性价比相对来说要不算最好 中规中矩 总的来说推荐购买。【其它描述】没有ESP和自动落锁 后排座椅不能放倒......不能再多说了 毕竟才10万的合资车。【为什么最终选择这款车】对比了昂克赛拉 起亚k3|朗动 轩逸 蓝鸟 朗逸这几款后 韩系车技术老旧被朋友给排除了；昂克赛拉虽然外观时尚 有创驰蓝天技术 但是自动挡要比卡罗拉贵2万 养护费用可能比卡罗拉要高 排除；轩逸和蓝鸟外配置相当 但新车没有啥优惠 排除；朗逸外观跟捷达一样 排除。最后在丰田故障率小 维护保养省钱 保值率高的口碑参考下选择了小卡。"|http://k.autohome.com.cn/spec/18890/view_1170228_1.html?st=104&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522345609|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 10:23:13|2016年06月26日 发表了口碑|来自：汽车之家iPhone版  2016年06月26日 发表了口碑  口碑   《卡罗拉的外观是我最看好的 当时再k3和卡罗拉做选选择》           【最满意的一点】手动档的车提速快 我喜欢提速的感觉 犀利的大灯 真是让人喜欢的不得了 我买的是外白内黑的 当时有一辆外白内黄的自动档的 我却没要【最不满意的一点】后来买完车交往了个女朋友 谁知媳妇的车是2011款马六 如果用两个车太浪费 她的怎么说也年岁久了 卖她那一部 可是我这个却是手动挡的 她说开着太费脑子 让现在的自动档气死了 以后大家谨记千万自动档 要不会有后悔的那天 开手动挡的 看着档次低【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】没有太中意的 直接看好这车了 直接去的莱州安利捷4s店【其他描述】|http://k.autohome.com.cn/spec/18891/view_1184866_1.html?st=3&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522443497|Autohome_review|뉴 보라(宝来)|ZHO|2016-06-27 11:25:19|2016年06月23日 发表了口碑|来自：手机汽车之家  2016年06月23日 发表了口碑  口碑   《稳固的德国工艺制作的底盘让弯道和颠簸路面不再那么困扰你。》   【最满意的一点】一般的油耗可以感受到大扭矩的动力。【最不满意的一点】内饰和外观设计中规中矩 想改装的部件较少。【空间】空间差异有点不足 宝来的价格桑塔纳的空间。【动力】动力杠杠的！宝来的价格近于高尔夫gti的享受【操控】前独立悬挂后连横式设计也是常规配置。【油耗】跟日系车没法比 相当于日系车安全性能也比不了一样。【舒适性】车内隔音效果相对比较不错的 【外观】个人比较喜欢外观改装的车型 宝来中规中矩外观改装的局限性很大。【内饰】座椅是高级仿pu的abs混合皮具 防龟裂较好 就是空间太不理想 宝来的价格桑塔纳的空间！【性价比】 总体来说宝来在同级车车里性价比很好 日系的卡罗拉ex 飞度 思域除了油耗低其他都是纸 韩系的k3 索纳塔 都是得个壳 国产的就不说了十几万买个国产仿制车没意思 法国和通用车那不是烧油是喝油。其他个各花入各眼【为什么最终选择这款车？】同价位的车对比中性价比很高 比国产 日 韩系车坚稳 比美国车省油。【其他描述】|http://k.autohome.com.cn/spec/14422/view_1181439_1.html?st=14&piap=0 633 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522524549|Autohome_review|닛산 티아나(天籁)|ZHO|2016-06-27 12:07:14|2016年06月20日 发表了口碑|来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《性价比超高 外观大气稳重 省油。》             【最满意的一点】坐椅舒适 减震不错 空间宽敞 电动坐椅 后排出风口非常好。【最不满意的一点】自动大反应慢 基本没用 舒适版无倒车雷达 好歹十几万的车 居然不配这个两百块钱又非常实用的东西？前保险杠与叶子板接合处是水平状态 下雨天开车后污垢会从接合处流到保险杠上 很难看 我观察过其他车 其他车的这个部位一般都是有一个角度的 污水会顺着角度流到地上 不会弄脏保险杠 我认为这是设计不到位。【空间】很满意 现在看别人家的车都觉得小【动力】比原来的1.4强多了。【操控】没开过其他车 反正比k2好【油耗】没k2省 不过排量大0.6车重四百公斤 很不错了。我最低开过3.6升百公里 一般来说两百块跑四百三四十公里 高速城区农村各有一部分 如果纯城区只能跑三百六十左右。【舒适性】不错 买天籁就是冲这个来的 我腰椎间盘突出 做了手术 上了钢筋的 不能受冲击 过减速带比原来好多了【外观】大气稳重【内饰】还行 有味 但比原车好。【性价比】超高 别人都说这车得二十几万吧 我说十五万没人信。【为什么最终选择这款车？】由于前一个车是起亚k2 所以最先看的是k3 媳妇试坐之后认为除了大点之外和k2没啥区别 后来又试了一些其他车 都没感觉 直到走进一家店里看到天籁 媳妇坐进去试了一下 感觉很满意 移沙发确实不错 但是就是觉得价格超了 那是去年的事了 今年三月又去试了kx3 板车悬挂同样让人不满意 本地车展又去转了转 带媳妇去看了丰田卡罗拉 内饰丑死个人 比老款难看多了 后来媳妇发话 干脆一步到位 上天籁。【其他描述】|http://k.autohome.com.cn/spec/15104/view_1173431_1.html?st=49&piap=0 634 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522545336|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 12:21:14|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=161&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522545465|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 12:21:14|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=147&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522545661|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 12:21:15|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=125&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522546142|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 12:21:24|2016年06月19日 发表了口碑|来自：手机汽车之家  2016年06月19日 发表了口碑  口碑    《外观好看.性价比不错》             【最满意的一点】动力可以.颜值不错.空间杠杠的！油耗在接受范围内……不到五毛一公里.【最不满意的一点】避震较硬..隔音不太好..换档不是太顺..还有最重要的一点这款车居然只有一条智能钥匙.起亚有点抠哦！【空间】空间杠杠的.驾驶位我一米七的身高座的好宽松 特别是后座中间凸起几乎可以忽略 比帝豪强多了 帝豪后面凸起真心好高。【动力】对于在城里跑动力真心够用 如果不在乎油耗的话 只要舍得踩油门动力要多少是多少。【操控】指向没什么问题 就是方向盘有点重 换挡时有点卡 倒车时好容易熄火。六档位开起来好爽！【油耗】加了200跑了460多公里 算下来不到五毛一公里。油耗还是可以的 只是论坛里他们开出3～4毛一公里.所以觉得我的油耗还是下降空间滴！【舒适性】座椅还可以 就是隔音不是很好【外观】满分 开卡罗拉的朋友说我这张好有宽体轿跑的感觉??????【内饰】塑料感有点强【性价比】性价比没的说！非常可以！特别是15款！【为什么最终选择这款车？】最初是看上哈佛h5的 .奈何钱包米不够再加上我们当地的哈佛4s店服务真的太差了.直接是鼻子登天牛B哄哄的（昆明迪鑫）以后我还会买哈佛但绝对不在这家店买！不好意思情不自禁偏题了????言归正传 后来又去看远景看着看着就帝豪.看完后都决定上帝豪了.就在去订车的途中朋友说起他们店的15款k3在搞活动算下来跟帝豪差不多价格.然后就掉头直奔起亚家.直到定了车我才去论坛了解这款车.还好论坛里都说这张车不错【其他描述】把小三带回家绝不后悔 你值得拥有！导航和真皮座椅都是提车后在外面做的。|http://k.autohome.com.cn/spec/19723/view_1172428_1.html?st=63&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522546197|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 12:21:24|2016年06月20日 发表了口碑|来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《前脸16新款看上去比15款锐利了…》             【最满意的一点】最满意的就是性价比了…优惠过后同样的配置价格低…【最不满意的一点】提速有点慢…每次等红灯 都要深踩油门  中控丑 后备箱垫子塌陷…问4s怎么解决 竟然告诉我东西放两边 不要放中间 好吧 你赢了…【空间】对空间比较满意…媳妇说后排比她妹妹家索八小不多少…【动力】动力给4分吧 毕竟排量小…不过也够用了 【操控】没开过太多车 不懂操控 不过已经很满足了 操控比两轮电动车爽 哈哈…??【油耗】还在磨合期 上了高速匀速80 最低油耗5.2 比较满意吧【舒适性】前排舒适度不错…大儿子把后排当沙发蹦来蹦去…由此可见后面还是不错 【外观】这个要给满分 外表很漂亮 个人感觉比15款好看…【内饰】内饰只能给3分…虽然说看习惯了 但还是想说一句：太丑了…【性价比】性价比无敌…16增加了ESP 10.6万的车送了导航皮座椅贴膜脚垫…空间大 配置高 价格合适…总体来说还是瑕不掩瑜的…【为什么最终选择这款车？】选车历程比较艰辛…两个儿子了 用钱的地方太多 只有精打细算 虽然很想支持国产 但第一辆车还是打算耐用点 日系卡罗拉 1.6竟然没有ESP 而且价格偏高 美系新英朗 因为没买车之前用车都是借的表哥英朗 油耗有点高 也不想买同一个车了 别的就不说了 反正各种原因pass掉了 关注起亚其实是看中kx3了 无奈价格有点接受不了 前一段表妹家提了k3 感觉还不错 就把目光转投k3 事实证明车还是很不错的…【其他描述】喜欢就下手吧 普遍优惠都在1.5万左右 …不会让你失望的|http://k.autohome.com.cn/spec/25739/view_1174824_1.html?st=53&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522564325|Autohome_review|포커스(福克斯)|ZHO|2016-06-27 12:30:04|2016年06月20日 发表了口碑|"来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《唯一缺点就是空间小！》           【最满意的一点】好开 很稳 很省心 【最不满意的一点】空间小 降价快【空间】坐五个人不是太挤 后备箱比较大 综合还是不错【动力】不开空调 一个人开还是不错的 要舍得给油！驾驶乐趣不错 满座来空调那就力不从心了【操控】转向精准 悬架支撑不错 过弯比较有信心 过坑洼路面不是太舒服！【油耗】油耗还能接受 不是太高！当然没发和日系车比咯！【舒适性】座椅包裹性好 不过长途驾驶感觉不太舒服 座椅不是太软。关窗静音效果不错 胎噪有点大 其他方面都还不错的！【外观】外观还是比较漂亮的！轮毂再大一号就帅多了！【内饰】用料不错 做工就不敢恭维了！缝隙太大 不像合资的车。哎！真是应征了网友们所说的?百年福特毁于长安！希望长安福特之后们在做工方面改善改善！【性价比】性能不错 安全配置比较齐全 长安的价格贬值比较快！很让消费者伤心??买了车快两年了 唯一后悔的就是不该买最低配版的 如果再给我重新选择的机会 毫不犹豫直接上中高配！！！！！！！！！！【为什么最终选择这款车？】朗动 k3|朗逸。朗动挺漂亮 老婆看的时候说感觉太单薄.k3和朗动差不懂 配置也差不多 朋友的也是k3|不想大家都买一样的 果断放弃。朗逸神车 比较中庸 保值率高 不适合我们九零后 要有个性。福克斯基本安全配置比较高 油耗必上一代有所改善 车身扎实。比较适合自己 空间勉强够用 主要是自己开 能接受。【其他描述】油箱负压 空调效果不是很好 保养贵"|http://k.autohome.com.cn/spec/12132/view_1176643_1.html?st=107&piap=0 364 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522597199|Autohome_review|닛산 티아나(天籁)|ZHO|2016-06-27 12:49:02|2016年06月20日 发表了口碑|来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《性价比超高 外观大气稳重 省油。》             【最满意的一点】坐椅舒适 减震不错 空间宽敞 电动坐椅 后排出风口非常好。【最不满意的一点】自动大反应慢 基本没用 舒适版无倒车雷达 好歹十几万的车 居然不配这个两百块钱又非常实用的东西？前保险杠与叶子板接合处是水平状态 下雨天开车后污垢会从接合处流到保险杠上 很难看 我观察过其他车 其他车的这个部位一般都是有一个角度的 污水会顺着角度流到地上 不会弄脏保险杠 我认为这是设计不到位。【空间】很满意 现在看别人家的车都觉得小【动力】比原来的1.4强多了。【操控】没开过其他车 反正比k2好【油耗】没k2省 不过排量大0.6车重四百公斤 很不错了。我最低开过3.6升百公里 一般来说两百块跑四百三四十公里 高速城区农村各有一部分 如果纯城区只能跑三百六十左右。【舒适性】不错 买天籁就是冲这个来的 我腰椎间盘突出 做了手术 上了钢筋的 不能受冲击 过减速带比原来好多了【外观】大气稳重【内饰】还行 有味 但比原车好。【性价比】超高 别人都说这车得二十几万吧 我说十五万没人信。【为什么最终选择这款车？】由于前一个车是起亚k2 所以最先看的是k3 媳妇试坐之后认为除了大点之外和k2没啥区别 后来又试了一些其他车 都没感觉 直到走进一家店里看到天籁 媳妇坐进去试了一下 感觉很满意 移沙发确实不错 但是就是觉得价格超了 那是去年的事了 今年三月又去试了kx3 板车悬挂同样让人不满意 本地车展又去转了转 带媳妇去看了丰田卡罗拉 内饰丑死个人 比老款难看多了 后来媳妇发话 干脆一步到位 上天籁。【其他描述】|http://k.autohome.com.cn/spec/15104/view_1173431_1.html?st=51&piap=0 634 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522617840|Autohome_review|포커스(福克斯)|ZHO|2016-06-27 13:03:04|2016年06月20日 发表了口碑|"来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《唯一缺点就是空间小！》           【最满意的一点】好开 很稳 很省心 【最不满意的一点】空间小 降价快【空间】坐五个人不是太挤 后备箱比较大 综合还是不错【动力】不开空调 一个人开还是不错的 要舍得给油！驾驶乐趣不错 满座来空调那就力不从心了【操控】转向精准 悬架支撑不错 过弯比较有信心 过坑洼路面不是太舒服！【油耗】油耗还能接受 不是太高！当然没发和日系车比咯！【舒适性】座椅包裹性好 不过长途驾驶感觉不太舒服 座椅不是太软。关窗静音效果不错 胎噪有点大 其他方面都还不错的！【外观】外观还是比较漂亮的！轮毂再大一号就帅多了！【内饰】用料不错 做工就不敢恭维了！缝隙太大 不像合资的车。哎！真是应征了网友们所说的?百年福特毁于长安！希望长安福特之后们在做工方面改善改善！【性价比】性能不错 安全配置比较齐全 长安的价格贬值比较快！很让消费者伤心??买了车快两年了 唯一后悔的就是不该买最低配版的 如果再给我重新选择的机会 毫不犹豫直接上中高配！！！！！！！！！！【为什么最终选择这款车？】朗动 k3|朗逸。朗动挺漂亮 老婆看的时候说感觉太单薄.k3和朗动差不懂 配置也差不多 朋友的也是k3|不想大家都买一样的 果断放弃。朗逸神车 比较中庸 保值率高 不适合我们九零后 要有个性。福克斯基本安全配置比较高 油耗必上一代有所改善 车身扎实。比较适合自己 空间勉强够用 主要是自己开 能接受。【其他描述】油箱负压 空调效果不是很好 保养贵"|http://k.autohome.com.cn/spec/12132/view_1176643_1.html?st=108&piap=0 364 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522649062|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 13:23:01|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=162&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522649076|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 13:23:01|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=148&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522649098|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 13:23:01|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=126&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522649162|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 13:23:01|2016年06月19日 发表了口碑|来自：手机汽车之家  2016年06月19日 发表了口碑  口碑    《外观好看.性价比不错》             【最满意的一点】动力可以.颜值不错.空间杠杠的！油耗在接受范围内……不到五毛一公里.【最不满意的一点】避震较硬..隔音不太好..换档不是太顺..还有最重要的一点这款车居然只有一条智能钥匙.起亚有点抠哦！【空间】空间杠杠的.驾驶位我一米七的身高座的好宽松 特别是后座中间凸起几乎可以忽略 比帝豪强多了 帝豪后面凸起真心好高。【动力】对于在城里跑动力真心够用 如果不在乎油耗的话 只要舍得踩油门动力要多少是多少。【操控】指向没什么问题 就是方向盘有点重 换挡时有点卡 倒车时好容易熄火。六档位开起来好爽！【油耗】加了200跑了460多公里 算下来不到五毛一公里。油耗还是可以的 只是论坛里他们开出3～4毛一公里.所以觉得我的油耗还是下降空间滴！【舒适性】座椅还可以 就是隔音不是很好【外观】满分 开卡罗拉的朋友说我这张好有宽体轿跑的感觉??????【内饰】塑料感有点强【性价比】性价比没的说！非常可以！特别是15款！【为什么最终选择这款车？】最初是看上哈佛h5的 .奈何钱包米不够再加上我们当地的哈佛4s店服务真的太差了.直接是鼻子登天牛B哄哄的（昆明迪鑫）以后我还会买哈佛但绝对不在这家店买！不好意思情不自禁偏题了????言归正传 后来又去看远景看着看着就帝豪.看完后都决定上帝豪了.就在去订车的途中朋友说起他们店的15款k3在搞活动算下来跟帝豪差不多价格.然后就掉头直奔起亚家.直到定了车我才去论坛了解这款车.还好论坛里都说这张车不错【其他描述】把小三带回家绝不后悔 你值得拥有！导航和真皮座椅都是提车后在外面做的。|http://k.autohome.com.cn/spec/19723/view_1172428_1.html?st=64&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522649172|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 13:23:01|2016年06月20日 发表了口碑|来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《前脸16新款看上去比15款锐利了…》             【最满意的一点】最满意的就是性价比了…优惠过后同样的配置价格低…【最不满意的一点】提速有点慢…每次等红灯 都要深踩油门  中控丑 后备箱垫子塌陷…问4s怎么解决 竟然告诉我东西放两边 不要放中间 好吧 你赢了…【空间】对空间比较满意…媳妇说后排比她妹妹家索八小不多少…【动力】动力给4分吧 毕竟排量小…不过也够用了 【操控】没开过太多车 不懂操控 不过已经很满足了 操控比两轮电动车爽 哈哈…??【油耗】还在磨合期 上了高速匀速80 最低油耗5.2 比较满意吧【舒适性】前排舒适度不错…大儿子把后排当沙发蹦来蹦去…由此可见后面还是不错 【外观】这个要给满分 外表很漂亮 个人感觉比15款好看…【内饰】内饰只能给3分…虽然说看习惯了 但还是想说一句：太丑了…【性价比】性价比无敌…16增加了ESP 10.6万的车送了导航皮座椅贴膜脚垫…空间大 配置高 价格合适…总体来说还是瑕不掩瑜的…【为什么最终选择这款车？】选车历程比较艰辛…两个儿子了 用钱的地方太多 只有精打细算 虽然很想支持国产 但第一辆车还是打算耐用点 日系卡罗拉 1.6竟然没有ESP 而且价格偏高 美系新英朗 因为没买车之前用车都是借的表哥英朗 油耗有点高 也不想买同一个车了 别的就不说了 反正各种原因pass掉了 关注起亚其实是看中kx3了 无奈价格有点接受不了 前一段表妹家提了k3 感觉还不错 就把目光转投k3 事实证明车还是很不错的…【其他描述】喜欢就下手吧 普遍优惠都在1.5万左右 …不会让你失望的|http://k.autohome.com.cn/spec/25739/view_1174824_1.html?st=54&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522706558|Autohome_review|랑동(朗动)|ZHO|2016-06-27 13:59:02|2016年06月21日 发表了口碑|来自：手机汽车之家  2016年06月21日 发表了口碑  口碑   《外观时尚好看 车子配置高实惠》           【最满意的一点】车子的外观和空间【最不满意的一点】1.6发动机动力不足【空间】后排虽然不能放倒 但足够日常生活所用 如何是放大东西的话就放不进去了【动力】起步肉 加速平稳 如果跑高速的话 油门响应有点慢 比如在跑高速过程中 你松下油门再想加速踩油门要踩深一点 中间有2秒的停顿加速【操控】方向盘轻 方向比较准【油耗】综合油耗还可以接受【舒适性】座椅很舒服 胎噪比较大跑高速【外观】外观非常喜欢【内饰】内饰中控台是软的比思域硬胶好很多【性价比】配置高 价格便宜实惠【为什么最终选择这款车？】选车中看了思域 速腾 卡罗拉 雷凌 k3。朗动的外观内饰价格优惠吸引我【其他描述】|http://k.autohome.com.cn/spec/20618/view_1178572_1.html?st=35&piap=0 2764 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522714605|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 14:05:01|2016年06月18日 发表了口碑|"2016年06月18日 发表了口碑  口碑    《空间大 省油 外观大气 优惠力度大》             【最满意的一点】空间大 油耗低 外观时尚 1万公里换机油保养。【最不满意的一点】没有ESP 没有发动机防盗 这俩项确实不应该简配。【空间】买车前参考过昂克赛拉 起亚k3|朗动 轩逸 蓝鸟 朗逸。轴距都是2700mm|但是看罗拉空间明显要大一些。180的大长腿坐进去都不挤。后排地面中间平整 也没有扶手 座三个175的壮汉也不觉得挤 不过后备箱不如轩逸的 感觉略小。【动力】1.6L的动力一个人开经常会有推背感 毕竟122马力 哈哈 但是座人了就感觉肉了 不过比朋友的斯柯达明锐1.6L双离合还是强劲不少 而且自然吸气的发动机跟涡轮增压比起来也没有烧机油的风险。【操控】之前开过面包车 开过荣威 但是跟卡罗拉的CVT比起来差远了 卡罗拉的标定确实比较扎实 换挡逻辑非常清新 开起来很平顺 出乎意料。在市区基本在1000转左右 处于ECO模式 高速跑120迈也就不到2000转左右 不知道需不需要像有的老司机说的过了磨合期高速拉缸。【油耗】刚提车时候油耗归零 开了110公里 竟然达到了惊人的4.1L/百公里 后来随着里程的增加逐步稳定在了6.5 6.6。日系车省油的名号确实不是盖的。【舒适性】这个价位的卡罗拉没有独立悬挂确实有些遗憾 在过减速带的时候 感觉略硬 风噪没有群友说的夸张 到了100迈内部还是比较安静的 但是偶尔能听到像石子刮地的声音 一直找不到原因。【外观】外观比老款的确实好看 个人觉得比雷凌的要收敛 离地间隙很低 好看但是也容易被磕碰。【内饰】内饰是硬塑料 黑白小仪表。10寸导航很加分 很大气 堪比K3.织物座椅去淘宝配个坐垫 美观舒适 朋友的真皮座椅夏天烫屁股。置物空间很多 放置杂物什么的没问题。【性价比】恰逢五一车展搞活动 优惠力度还是比较大了 送了贴膜导航装具行车记录仪。性价比相对来说要不算最好 中规中矩 总的来说推荐购买。【其它描述】没有ESP和自动落锁 后排座椅不能放倒......不能再多说了 毕竟才10万的合资车。【为什么最终选择这款车】对比了昂克赛拉 起亚k3|朗动 轩逸 蓝鸟 朗逸这几款后 韩系车技术老旧被朋友给排除了；昂克赛拉虽然外观时尚 有创驰蓝天技术 但是自动挡要比卡罗拉贵2万 养护费用可能比卡罗拉要高 排除；轩逸和蓝鸟外配置相当 但新车没有啥优惠 排除；朗逸外观跟捷达一样 排除。最后在丰田故障率小 维护保养省钱 保值率高的口碑参考下选择了小卡。"|http://k.autohome.com.cn/spec/18890/view_1170228_1.html?st=106&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522714721|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 14:05:02|2016年06月26日 发表了口碑|来自：汽车之家iPhone版  2016年06月26日 发表了口碑  口碑   《卡罗拉的外观是我最看好的 当时再k3和卡罗拉做选选择》           【最满意的一点】手动档的车提速快 我喜欢提速的感觉 犀利的大灯 真是让人喜欢的不得了 我买的是外白内黑的 当时有一辆外白内黄的自动档的 我却没要【最不满意的一点】后来买完车交往了个女朋友 谁知媳妇的车是2011款马六 如果用两个车太浪费 她的怎么说也年岁久了 卖她那一部 可是我这个却是手动挡的 她说开着太费脑子 让现在的自动档气死了 以后大家谨记千万自动档 要不会有后悔的那天 开手动挡的 看着档次低【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】没有太中意的 直接看好这车了 直接去的莱州安利捷4s店【其他描述】|http://k.autohome.com.cn/spec/18891/view_1184866_1.html?st=5&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522761967|Autohome_review|포커스(福克斯)|ZHO|2016-06-27 14:32:02|2016年06月20日 发表了口碑|"来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《唯一缺点就是空间小！》           【最满意的一点】好开 很稳 很省心 【最不满意的一点】空间小 降价快【空间】坐五个人不是太挤 后备箱比较大 综合还是不错【动力】不开空调 一个人开还是不错的 要舍得给油！驾驶乐趣不错 满座来空调那就力不从心了【操控】转向精准 悬架支撑不错 过弯比较有信心 过坑洼路面不是太舒服！【油耗】油耗还能接受 不是太高！当然没发和日系车比咯！【舒适性】座椅包裹性好 不过长途驾驶感觉不太舒服 座椅不是太软。关窗静音效果不错 胎噪有点大 其他方面都还不错的！【外观】外观还是比较漂亮的！轮毂再大一号就帅多了！【内饰】用料不错 做工就不敢恭维了！缝隙太大 不像合资的车。哎！真是应征了网友们所说的?百年福特毁于长安！希望长安福特之后们在做工方面改善改善！【性价比】性能不错 安全配置比较齐全 长安的价格贬值比较快！很让消费者伤心??买了车快两年了 唯一后悔的就是不该买最低配版的 如果再给我重新选择的机会 毫不犹豫直接上中高配！！！！！！！！！！【为什么最终选择这款车？】朗动 k3|朗逸。朗动挺漂亮 老婆看的时候说感觉太单薄.k3和朗动差不懂 配置也差不多 朋友的也是k3|不想大家都买一样的 果断放弃。朗逸神车 比较中庸 保值率高 不适合我们九零后 要有个性。福克斯基本安全配置比较高 油耗必上一代有所改善 车身扎实。比较适合自己 空间勉强够用 主要是自己开 能接受。【其他描述】油箱负压 空调效果不是很好 保养贵"|http://k.autohome.com.cn/spec/12132/view_1176643_1.html?st=109&piap=0 364 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522782857|Autohome_review|아반떼 AD(领动)|ZHO|2016-06-27 14:44:03|2016年06月02日 发表了口碑|来自：手机汽车之家  2016年06月02日 发表了口碑  口碑    《外观拉风 配置足够 整体性价比还是不错的。》           【最满意的一点】外观很拉风 现在路上还很少见 大轮毂。日间行车灯很高大上 自动头灯也很高端。中控台是软的 车内显示屏清晰度很高。倒车影像有随动辅助导线。很方便。车内音响很赞 我喜欢听音乐 完全满足我的要求。【最不满意的一点】后排不能放倒 这个真心很郁闷 这个放倒真的很难吗？这几天B柱内有异响 这还是新车呀 哎。。过几天去4s看看 希望不是啥大问题。另外胎噪确实大 我想跟轮胎大也有关系吧。悬挂还是有点硬 不过在接受范围内。【空间】空间同级别还是有优势的 中间无凸起。【动力】动力够用 现在用的eco模式【操控】转向精准 没啥虚位。【油耗】表显6 肯定是不准的 等下次油表亮再算算。【舒适性】还可以 家用够了。【外观】满意【内饰】做工还是比较好的 接缝均匀。【性价比】性价比高【为什么最终选择这款车？】同级别都看了 也试驾了 福克斯空间太小 科鲁兹都说油耗高 新英朗有点老气 卡罗拉没esp 思域根本没现车 看来看去家用也就韩系车了。【其他描述】换车的想法去年就有了 但是一直没有付诸行动 一是因为暂时有车开 二是今年上市新车多 想再等等 经常看论坛 心里已经有了几个备选 英朗 老表刚买的 开始觉得性价比很高 后来发现新旧差别很大 就pass了。福克斯外观不错 但是同事有好几辆 不想买一样的。k3性价比很高 优惠很大 但是新款感觉你没老款好看。看到最后就是领动了 配置高 外观拉风 总体性价比很高。|http://k.autohome.com.cn/spec/25701/view_1148059_1.html?st=112&piap=0 3959 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522783004|Autohome_review|아반떼 AD(领动)|ZHO|2016-06-27 14:44:04|2016年06月19日 发表了口碑|来自：手机汽车之家  2016年06月19日 发表了口碑  口碑    《选择不后悔 领动 领新而动。》             【最满意的一点】配置够用 外观造型动感。油耗表现好。磨合期过了后应该到正常水平了 现在降到8.3L了。【最不满意的一点】暂时还没发现 非要说的话速度上来后有点胎噪 另外轮胎有点卡小石子。【空间】我觉得空间很大了 后排的同事说不压抑 空间宽敞。头部空间和腿部空间都很充足 我身高173cm 不错。【动力】动力充足 只要肯给油 深踩油门 立马就走 反应灵敏 还没体验过运动模式 等磨合期完了试试。试驾的时候销售用1.4T的运动模式开过 感觉动力很猛。【操控】转向系统反应灵敏 方向盘虚位少 指向精准。悬架系统支撑性好 很稳。我在试驾的时候销售特地带我体验了一下转急弯 没有一点多余的倾斜。【油耗】刚提车的时候是18.几 慢慢的降下来了。满足预期 目前在磨合期 油耗下来了。【舒适性】座椅挺舒服的 我没加装真皮 感觉够用了。【外观】外观拉风 特别是前脸造型。【内饰】内饰设计很用心 能够平常接触的地方都是软材料 用心去体验啦。【性价比】自动精英版本配置够用了 具体的可以去看参数 选择不后悔。目前虽然没有大的降价 但是早买早享受了。【为什么最终选择这款车？】一直纠结着到底买哪款 去4s店看了好多车型 选车的时候看了卡罗拉 雷凌 起亚k3 领动 朗动 最终选择了领动 新款 1.6L购置税减半 自动精英型配置够用了。满意。另外就是感觉领动挺符合年轻人的气质的。我今年26岁 感觉其他车型不太符合 有的太中庸 有的太成熟了。这个刚刚好。还有就是胡歌代言的 挺喜欢胡歌的 哈哈 花痴了。【其他描述】今天看到了2辆白色的领动 对了 我定车那天4s店里的一台展车柠檬黄被人买了 很拉风。|http://k.autohome.com.cn/spec/25701/view_1171797_1.html?st=56&piap=0 3959 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522795455|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 14:52:02|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=164&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522795490|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 14:52:02|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=150&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522795546|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 14:52:02|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=128&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522795700|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 14:52:02|2016年06月19日 发表了口碑|来自：手机汽车之家  2016年06月19日 发表了口碑  口碑    《外观好看.性价比不错》             【最满意的一点】动力可以.颜值不错.空间杠杠的！油耗在接受范围内……不到五毛一公里.【最不满意的一点】避震较硬..隔音不太好..换档不是太顺..还有最重要的一点这款车居然只有一条智能钥匙.起亚有点抠哦！【空间】空间杠杠的.驾驶位我一米七的身高座的好宽松 特别是后座中间凸起几乎可以忽略 比帝豪强多了 帝豪后面凸起真心好高。【动力】对于在城里跑动力真心够用 如果不在乎油耗的话 只要舍得踩油门动力要多少是多少。【操控】指向没什么问题 就是方向盘有点重 换挡时有点卡 倒车时好容易熄火。六档位开起来好爽！【油耗】加了200跑了460多公里 算下来不到五毛一公里。油耗还是可以的 只是论坛里他们开出3～4毛一公里.所以觉得我的油耗还是下降空间滴！【舒适性】座椅还可以 就是隔音不是很好【外观】满分 开卡罗拉的朋友说我这张好有宽体轿跑的感觉??????【内饰】塑料感有点强【性价比】性价比没的说！非常可以！特别是15款！【为什么最终选择这款车？】最初是看上哈佛h5的 .奈何钱包米不够再加上我们当地的哈佛4s店服务真的太差了.直接是鼻子登天牛B哄哄的（昆明迪鑫）以后我还会买哈佛但绝对不在这家店买！不好意思情不自禁偏题了????言归正传 后来又去看远景看着看着就帝豪.看完后都决定上帝豪了.就在去订车的途中朋友说起他们店的15款k3在搞活动算下来跟帝豪差不多价格.然后就掉头直奔起亚家.直到定了车我才去论坛了解这款车.还好论坛里都说这张车不错【其他描述】把小三带回家绝不后悔 你值得拥有！导航和真皮座椅都是提车后在外面做的。|http://k.autohome.com.cn/spec/19723/view_1172428_1.html?st=66&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522795726|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 14:52:02|2016年06月20日 发表了口碑|来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《前脸16新款看上去比15款锐利了…》             【最满意的一点】最满意的就是性价比了…优惠过后同样的配置价格低…【最不满意的一点】提速有点慢…每次等红灯 都要深踩油门  中控丑 后备箱垫子塌陷…问4s怎么解决 竟然告诉我东西放两边 不要放中间 好吧 你赢了…【空间】对空间比较满意…媳妇说后排比她妹妹家索八小不多少…【动力】动力给4分吧 毕竟排量小…不过也够用了 【操控】没开过太多车 不懂操控 不过已经很满足了 操控比两轮电动车爽 哈哈…??【油耗】还在磨合期 上了高速匀速80 最低油耗5.2 比较满意吧【舒适性】前排舒适度不错…大儿子把后排当沙发蹦来蹦去…由此可见后面还是不错 【外观】这个要给满分 外表很漂亮 个人感觉比15款好看…【内饰】内饰只能给3分…虽然说看习惯了 但还是想说一句：太丑了…【性价比】性价比无敌…16增加了ESP 10.6万的车送了导航皮座椅贴膜脚垫…空间大 配置高 价格合适…总体来说还是瑕不掩瑜的…【为什么最终选择这款车？】选车历程比较艰辛…两个儿子了 用钱的地方太多 只有精打细算 虽然很想支持国产 但第一辆车还是打算耐用点 日系卡罗拉 1.6竟然没有ESP 而且价格偏高 美系新英朗 因为没买车之前用车都是借的表哥英朗 油耗有点高 也不想买同一个车了 别的就不说了 反正各种原因pass掉了 关注起亚其实是看中kx3了 无奈价格有点接受不了 前一段表妹家提了k3 感觉还不错 就把目光转投k3 事实证明车还是很不错的…【其他描述】喜欢就下手吧 普遍优惠都在1.5万左右 …不会让你失望的|http://k.autohome.com.cn/spec/25739/view_1174824_1.html?st=56&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522805383|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 14:57:03|2016年06月18日 发表了口碑|"2016年06月18日 发表了口碑  口碑    《空间大 省油 外观大气 优惠力度大》             【最满意的一点】空间大 油耗低 外观时尚 1万公里换机油保养。【最不满意的一点】没有ESP 没有发动机防盗 这俩项确实不应该简配。【空间】买车前参考过昂克赛拉 起亚k3|朗动 轩逸 蓝鸟 朗逸。轴距都是2700mm|但是看罗拉空间明显要大一些。180的大长腿坐进去都不挤。后排地面中间平整 也没有扶手 座三个175的壮汉也不觉得挤 不过后备箱不如轩逸的 感觉略小。【动力】1.6L的动力一个人开经常会有推背感 毕竟122马力 哈哈 但是座人了就感觉肉了 不过比朋友的斯柯达明锐1.6L双离合还是强劲不少 而且自然吸气的发动机跟涡轮增压比起来也没有烧机油的风险。【操控】之前开过面包车 开过荣威 但是跟卡罗拉的CVT比起来差远了 卡罗拉的标定确实比较扎实 换挡逻辑非常清新 开起来很平顺 出乎意料。在市区基本在1000转左右 处于ECO模式 高速跑120迈也就不到2000转左右 不知道需不需要像有的老司机说的过了磨合期高速拉缸。【油耗】刚提车时候油耗归零 开了110公里 竟然达到了惊人的4.1L/百公里 后来随着里程的增加逐步稳定在了6.5 6.6。日系车省油的名号确实不是盖的。【舒适性】这个价位的卡罗拉没有独立悬挂确实有些遗憾 在过减速带的时候 感觉略硬 风噪没有群友说的夸张 到了100迈内部还是比较安静的 但是偶尔能听到像石子刮地的声音 一直找不到原因。【外观】外观比老款的确实好看 个人觉得比雷凌的要收敛 离地间隙很低 好看但是也容易被磕碰。【内饰】内饰是硬塑料 黑白小仪表。10寸导航很加分 很大气 堪比K3.织物座椅去淘宝配个坐垫 美观舒适 朋友的真皮座椅夏天烫屁股。置物空间很多 放置杂物什么的没问题。【性价比】恰逢五一车展搞活动 优惠力度还是比较大了 送了贴膜导航装具行车记录仪。性价比相对来说要不算最好 中规中矩 总的来说推荐购买。【其它描述】没有ESP和自动落锁 后排座椅不能放倒......不能再多说了 毕竟才10万的合资车。【为什么最终选择这款车】对比了昂克赛拉 起亚k3|朗动 轩逸 蓝鸟 朗逸这几款后 韩系车技术老旧被朋友给排除了；昂克赛拉虽然外观时尚 有创驰蓝天技术 但是自动挡要比卡罗拉贵2万 养护费用可能比卡罗拉要高 排除；轩逸和蓝鸟外配置相当 但新车没有啥优惠 排除；朗逸外观跟捷达一样 排除。最后在丰田故障率小 维护保养省钱 保值率高的口碑参考下选择了小卡。"|http://k.autohome.com.cn/spec/18890/view_1170228_1.html?st=107&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522805645|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 14:57:04|2016年06月26日 发表了口碑|来自：汽车之家iPhone版  2016年06月26日 发表了口碑  口碑   《卡罗拉的外观是我最看好的 当时再k3和卡罗拉做选选择》           【最满意的一点】手动档的车提速快 我喜欢提速的感觉 犀利的大灯 真是让人喜欢的不得了 我买的是外白内黑的 当时有一辆外白内黄的自动档的 我却没要【最不满意的一点】后来买完车交往了个女朋友 谁知媳妇的车是2011款马六 如果用两个车太浪费 她的怎么说也年岁久了 卖她那一部 可是我这个却是手动挡的 她说开着太费脑子 让现在的自动档气死了 以后大家谨记千万自动档 要不会有后悔的那天 开手动挡的 看着档次低【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】没有太中意的 直接看好这车了 直接去的莱州安利捷4s店【其他描述】|http://k.autohome.com.cn/spec/18891/view_1184866_1.html?st=6&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522865414|Autohome_review|랑동(朗动)|ZHO|2016-06-27 15:32:02|2016年06月21日 发表了口碑|来自：手机汽车之家  2016年06月21日 发表了口碑  口碑   《外观时尚好看 车子配置高实惠》           【最满意的一点】车子的外观和空间【最不满意的一点】1.6发动机动力不足【空间】后排虽然不能放倒 但足够日常生活所用 如何是放大东西的话就放不进去了【动力】起步肉 加速平稳 如果跑高速的话 油门响应有点慢 比如在跑高速过程中 你松下油门再想加速踩油门要踩深一点 中间有2秒的停顿加速【操控】方向盘轻 方向比较准【油耗】综合油耗还可以接受【舒适性】座椅很舒服 胎噪比较大跑高速【外观】外观非常喜欢【内饰】内饰中控台是软的比思域硬胶好很多【性价比】配置高 价格便宜实惠【为什么最终选择这款车？】选车中看了思域 速腾 卡罗拉 雷凌 k3。朗动的外观内饰价格优惠吸引我【其他描述】|http://k.autohome.com.cn/spec/20618/view_1178572_1.html?st=36&piap=0 2764 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522877411|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 15:39:05|2016年06月18日 发表了口碑|"2016年06月18日 发表了口碑  口碑    《空间大 省油 外观大气 优惠力度大》             【最满意的一点】空间大 油耗低 外观时尚 1万公里换机油保养。【最不满意的一点】没有ESP 没有发动机防盗 这俩项确实不应该简配。【空间】买车前参考过昂克赛拉 起亚k3|朗动 轩逸 蓝鸟 朗逸。轴距都是2700mm|但是看罗拉空间明显要大一些。180的大长腿坐进去都不挤。后排地面中间平整 也没有扶手 座三个175的壮汉也不觉得挤 不过后备箱不如轩逸的 感觉略小。【动力】1.6L的动力一个人开经常会有推背感 毕竟122马力 哈哈 但是座人了就感觉肉了 不过比朋友的斯柯达明锐1.6L双离合还是强劲不少 而且自然吸气的发动机跟涡轮增压比起来也没有烧机油的风险。【操控】之前开过面包车 开过荣威 但是跟卡罗拉的CVT比起来差远了 卡罗拉的标定确实比较扎实 换挡逻辑非常清新 开起来很平顺 出乎意料。在市区基本在1000转左右 处于ECO模式 高速跑120迈也就不到2000转左右 不知道需不需要像有的老司机说的过了磨合期高速拉缸。【油耗】刚提车时候油耗归零 开了110公里 竟然达到了惊人的4.1L/百公里 后来随着里程的增加逐步稳定在了6.5 6.6。日系车省油的名号确实不是盖的。【舒适性】这个价位的卡罗拉没有独立悬挂确实有些遗憾 在过减速带的时候 感觉略硬 风噪没有群友说的夸张 到了100迈内部还是比较安静的 但是偶尔能听到像石子刮地的声音 一直找不到原因。【外观】外观比老款的确实好看 个人觉得比雷凌的要收敛 离地间隙很低 好看但是也容易被磕碰。【内饰】内饰是硬塑料 黑白小仪表。10寸导航很加分 很大气 堪比K3.织物座椅去淘宝配个坐垫 美观舒适 朋友的真皮座椅夏天烫屁股。置物空间很多 放置杂物什么的没问题。【性价比】恰逢五一车展搞活动 优惠力度还是比较大了 送了贴膜导航装具行车记录仪。性价比相对来说要不算最好 中规中矩 总的来说推荐购买。【其它描述】没有ESP和自动落锁 后排座椅不能放倒......不能再多说了 毕竟才10万的合资车。【为什么最终选择这款车】对比了昂克赛拉 起亚k3|朗动 轩逸 蓝鸟 朗逸这几款后 韩系车技术老旧被朋友给排除了；昂克赛拉虽然外观时尚 有创驰蓝天技术 但是自动挡要比卡罗拉贵2万 养护费用可能比卡罗拉要高 排除；轩逸和蓝鸟外配置相当 但新车没有啥优惠 排除；朗逸外观跟捷达一样 排除。最后在丰田故障率小 维护保养省钱 保值率高的口碑参考下选择了小卡。"|http://k.autohome.com.cn/spec/18890/view_1170228_1.html?st=108&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2522877690|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 15:39:05|2016年06月26日 发表了口碑|来自：汽车之家iPhone版  2016年06月26日 发表了口碑  口碑   《卡罗拉的外观是我最看好的 当时再k3和卡罗拉做选选择》           【最满意的一点】手动档的车提速快 我喜欢提速的感觉 犀利的大灯 真是让人喜欢的不得了 我买的是外白内黑的 当时有一辆外白内黄的自动档的 我却没要【最不满意的一点】后来买完车交往了个女朋友 谁知媳妇的车是2011款马六 如果用两个车太浪费 她的怎么说也年岁久了 卖她那一部 可是我这个却是手动挡的 她说开着太费脑子 让现在的自动档气死了 以后大家谨记千万自动档 要不会有后悔的那天 开手动挡的 看着档次低【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】没有太中意的 直接看好这车了 直接去的莱州安利捷4s店【其他描述】|http://k.autohome.com.cn/spec/18891/view_1184866_1.html?st=7&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523002741|Autohome_review|랑동(朗动)|ZHO|2016-06-27 16:48:04|2016年06月21日 发表了口碑|来自：手机汽车之家  2016年06月21日 发表了口碑  口碑   《外观时尚好看 车子配置高实惠》           【最满意的一点】车子的外观和空间【最不满意的一点】1.6发动机动力不足【空间】后排虽然不能放倒 但足够日常生活所用 如何是放大东西的话就放不进去了【动力】起步肉 加速平稳 如果跑高速的话 油门响应有点慢 比如在跑高速过程中 你松下油门再想加速踩油门要踩深一点 中间有2秒的停顿加速【操控】方向盘轻 方向比较准【油耗】综合油耗还可以接受【舒适性】座椅很舒服 胎噪比较大跑高速【外观】外观非常喜欢【内饰】内饰中控台是软的比思域硬胶好很多【性价比】配置高 价格便宜实惠【为什么最终选择这款车？】选车中看了思域 速腾 卡罗拉 雷凌 k3。朗动的外观内饰价格优惠吸引我【其他描述】|http://k.autohome.com.cn/spec/20618/view_1178572_1.html?st=37&piap=0 2764 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523020242|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 16:56:03|2016年06月26日 发表了口碑|来自：汽车之家iPhone版  2016年06月26日 发表了口碑  口碑   《卡罗拉的外观是我最看好的 当时再k3和卡罗拉做选选择》           【最满意的一点】手动档的车提速快 我喜欢提速的感觉 犀利的大灯 真是让人喜欢的不得了 我买的是外白内黑的 当时有一辆外白内黄的自动档的 我却没要【最不满意的一点】后来买完车交往了个女朋友 谁知媳妇的车是2011款马六 如果用两个车太浪费 她的怎么说也年岁久了 卖她那一部 可是我这个却是手动挡的 她说开着太费脑子 让现在的自动档气死了 以后大家谨记千万自动档 要不会有后悔的那天 开手动挡的 看着档次低【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】没有太中意的 直接看好这车了 直接去的莱州安利捷4s店【其他描述】|http://k.autohome.com.cn/spec/18891/view_1184866_1.html?st=8&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523026714|Autohome_review|뉴 보라(宝来)|ZHO|2016-06-27 17:00:01|2016年06月23日 发表了口碑|来自：手机汽车之家  2016年06月23日 发表了口碑  口碑   《稳固的德国工艺制作的底盘让弯道和颠簸路面不再那么困扰你。》   【最满意的一点】一般的油耗可以感受到大扭矩的动力。【最不满意的一点】内饰和外观设计中规中矩 想改装的部件较少。【空间】空间差异有点不足 宝来的价格桑塔纳的空间。【动力】动力杠杠的！宝来的价格近于高尔夫gti的享受【操控】前独立悬挂后连横式设计也是常规配置。【油耗】跟日系车没法比 相当于日系车安全性能也比不了一样。【舒适性】车内隔音效果相对比较不错的 【外观】个人比较喜欢外观改装的车型 宝来中规中矩外观改装的局限性很大。【内饰】座椅是高级仿pu的abs混合皮具 防龟裂较好 就是空间太不理想 宝来的价格桑塔纳的空间！【性价比】 总体来说宝来在同级车车里性价比很好 日系的卡罗拉ex 飞度 思域除了油耗低其他都是纸 韩系的k3 索纳塔 都是得个壳 国产的就不说了十几万买个国产仿制车没意思 法国和通用车那不是烧油是喝油。其他个各花入各眼【为什么最终选择这款车？】同价位的车对比中性价比很高 比国产 日 韩系车坚稳 比美国车省油。【其他描述】|http://k.autohome.com.cn/spec/14422/view_1181439_1.html?st=15&piap=0 633 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523038984|Autohome_review|포커스(福克斯)|ZHO|2016-06-27 17:07:35|2016年06月20日 发表了口碑|"来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《唯一缺点就是空间小！》           【最满意的一点】好开 很稳 很省心 【最不满意的一点】空间小 降价快【空间】坐五个人不是太挤 后备箱比较大 综合还是不错【动力】不开空调 一个人开还是不错的 要舍得给油！驾驶乐趣不错 满座来空调那就力不从心了【操控】转向精准 悬架支撑不错 过弯比较有信心 过坑洼路面不是太舒服！【油耗】油耗还能接受 不是太高！当然没发和日系车比咯！【舒适性】座椅包裹性好 不过长途驾驶感觉不太舒服 座椅不是太软。关窗静音效果不错 胎噪有点大 其他方面都还不错的！【外观】外观还是比较漂亮的！轮毂再大一号就帅多了！【内饰】用料不错 做工就不敢恭维了！缝隙太大 不像合资的车。哎！真是应征了网友们所说的?百年福特毁于长安！希望长安福特之后们在做工方面改善改善！【性价比】性能不错 安全配置比较齐全 长安的价格贬值比较快！很让消费者伤心??买了车快两年了 唯一后悔的就是不该买最低配版的 如果再给我重新选择的机会 毫不犹豫直接上中高配！！！！！！！！！！【为什么最终选择这款车？】朗动 k3|朗逸。朗动挺漂亮 老婆看的时候说感觉太单薄.k3和朗动差不懂 配置也差不多 朋友的也是k3|不想大家都买一样的 果断放弃。朗逸神车 比较中庸 保值率高 不适合我们九零后 要有个性。福克斯基本安全配置比较高 油耗必上一代有所改善 车身扎实。比较适合自己 空间勉强够用 主要是自己开 能接受。【其他描述】油箱负压 空调效果不是很好 保养贵"|http://k.autohome.com.cn/spec/12132/view_1176643_1.html?st=110&piap=0 364 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523095822|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 17:37:01|2016年06月26日 发表了口碑|来自：汽车之家iPhone版  2016年06月26日 发表了口碑  口碑   《卡罗拉的外观是我最看好的 当时再k3和卡罗拉做选选择》           【最满意的一点】手动档的车提速快 我喜欢提速的感觉 犀利的大灯 真是让人喜欢的不得了 我买的是外白内黑的 当时有一辆外白内黄的自动档的 我却没要【最不满意的一点】后来买完车交往了个女朋友 谁知媳妇的车是2011款马六 如果用两个车太浪费 她的怎么说也年岁久了 卖她那一部 可是我这个却是手动挡的 她说开着太费脑子 让现在的自动档气死了 以后大家谨记千万自动档 要不会有后悔的那天 开手动挡的 看着档次低【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】没有太中意的 直接看好这车了 直接去的莱州安利捷4s店【其他描述】|http://k.autohome.com.cn/spec/18891/view_1184866_1.html?st=9&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523146776|Autohome_review|닛산 티아나(天籁)|ZHO|2016-06-27 18:04:03|2016年06月20日 发表了口碑|来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《性价比超高 外观大气稳重 省油。》             【最满意的一点】坐椅舒适 减震不错 空间宽敞 电动坐椅 后排出风口非常好。【最不满意的一点】自动大反应慢 基本没用 舒适版无倒车雷达 好歹十几万的车 居然不配这个两百块钱又非常实用的东西？前保险杠与叶子板接合处是水平状态 下雨天开车后污垢会从接合处流到保险杠上 很难看 我观察过其他车 其他车的这个部位一般都是有一个角度的 污水会顺着角度流到地上 不会弄脏保险杠 我认为这是设计不到位。【空间】很满意 现在看别人家的车都觉得小【动力】比原来的1.4强多了。【操控】没开过其他车 反正比k2好【油耗】没k2省 不过排量大0.6车重四百公斤 很不错了。我最低开过3.6升百公里 一般来说两百块跑四百三四十公里 高速城区农村各有一部分 如果纯城区只能跑三百六十左右。【舒适性】不错 买天籁就是冲这个来的 我腰椎间盘突出 做了手术 上了钢筋的 不能受冲击 过减速带比原来好多了【外观】大气稳重【内饰】还行 有味 但比原车好。【性价比】超高 别人都说这车得二十几万吧 我说十五万没人信。【为什么最终选择这款车？】由于前一个车是起亚k2 所以最先看的是k3 媳妇试坐之后认为除了大点之外和k2没啥区别 后来又试了一些其他车 都没感觉 直到走进一家店里看到天籁 媳妇坐进去试了一下 感觉很满意 移沙发确实不错 但是就是觉得价格超了 那是去年的事了 今年三月又去试了kx3 板车悬挂同样让人不满意 本地车展又去转了转 带媳妇去看了丰田卡罗拉 内饰丑死个人 比老款难看多了 后来媳妇发话 干脆一步到位 上天籁。【其他描述】|http://k.autohome.com.cn/spec/15104/view_1173431_1.html?st=52&piap=0 634 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523168372|Autohome_review|포커스(福克斯)|ZHO|2016-06-27 18:17:53|2016年06月20日 发表了口碑|"来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《唯一缺点就是空间小！》           【最满意的一点】好开 很稳 很省心 【最不满意的一点】空间小 降价快【空间】坐五个人不是太挤 后备箱比较大 综合还是不错【动力】不开空调 一个人开还是不错的 要舍得给油！驾驶乐趣不错 满座来空调那就力不从心了【操控】转向精准 悬架支撑不错 过弯比较有信心 过坑洼路面不是太舒服！【油耗】油耗还能接受 不是太高！当然没发和日系车比咯！【舒适性】座椅包裹性好 不过长途驾驶感觉不太舒服 座椅不是太软。关窗静音效果不错 胎噪有点大 其他方面都还不错的！【外观】外观还是比较漂亮的！轮毂再大一号就帅多了！【内饰】用料不错 做工就不敢恭维了！缝隙太大 不像合资的车。哎！真是应征了网友们所说的?百年福特毁于长安！希望长安福特之后们在做工方面改善改善！【性价比】性能不错 安全配置比较齐全 长安的价格贬值比较快！很让消费者伤心??买了车快两年了 唯一后悔的就是不该买最低配版的 如果再给我重新选择的机会 毫不犹豫直接上中高配！！！！！！！！！！【为什么最终选择这款车？】朗动 k3|朗逸。朗动挺漂亮 老婆看的时候说感觉太单薄.k3和朗动差不懂 配置也差不多 朋友的也是k3|不想大家都买一样的 果断放弃。朗逸神车 比较中庸 保值率高 不适合我们九零后 要有个性。福克斯基本安全配置比较高 油耗必上一代有所改善 车身扎实。比较适合自己 空间勉强够用 主要是自己开 能接受。【其他描述】油箱负压 空调效果不是很好 保养贵"|http://k.autohome.com.cn/spec/12132/view_1176643_1.html?st=111&piap=0 364 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523174690|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 18:19:18|2016年06月18日 发表了口碑|"2016年06月18日 发表了口碑  口碑    《空间大 省油 外观大气 优惠力度大》             【最满意的一点】空间大 油耗低 外观时尚 1万公里换机油保养。【最不满意的一点】没有ESP 没有发动机防盗 这俩项确实不应该简配。【空间】买车前参考过昂克赛拉 起亚k3|朗动 轩逸 蓝鸟 朗逸。轴距都是2700mm|但是看罗拉空间明显要大一些。180的大长腿坐进去都不挤。后排地面中间平整 也没有扶手 座三个175的壮汉也不觉得挤 不过后备箱不如轩逸的 感觉略小。【动力】1.6L的动力一个人开经常会有推背感 毕竟122马力 哈哈 但是座人了就感觉肉了 不过比朋友的斯柯达明锐1.6L双离合还是强劲不少 而且自然吸气的发动机跟涡轮增压比起来也没有烧机油的风险。【操控】之前开过面包车 开过荣威 但是跟卡罗拉的CVT比起来差远了 卡罗拉的标定确实比较扎实 换挡逻辑非常清新 开起来很平顺 出乎意料。在市区基本在1000转左右 处于ECO模式 高速跑120迈也就不到2000转左右 不知道需不需要像有的老司机说的过了磨合期高速拉缸。【油耗】刚提车时候油耗归零 开了110公里 竟然达到了惊人的4.1L/百公里 后来随着里程的增加逐步稳定在了6.5 6.6。日系车省油的名号确实不是盖的。【舒适性】这个价位的卡罗拉没有独立悬挂确实有些遗憾 在过减速带的时候 感觉略硬 风噪没有群友说的夸张 到了100迈内部还是比较安静的 但是偶尔能听到像石子刮地的声音 一直找不到原因。【外观】外观比老款的确实好看 个人觉得比雷凌的要收敛 离地间隙很低 好看但是也容易被磕碰。【内饰】内饰是硬塑料 黑白小仪表。10寸导航很加分 很大气 堪比K3.织物座椅去淘宝配个坐垫 美观舒适 朋友的真皮座椅夏天烫屁股。置物空间很多 放置杂物什么的没问题。【性价比】恰逢五一车展搞活动 优惠力度还是比较大了 送了贴膜导航装具行车记录仪。性价比相对来说要不算最好 中规中矩 总的来说推荐购买。【其它描述】没有ESP和自动落锁 后排座椅不能放倒......不能再多说了 毕竟才10万的合资车。【为什么最终选择这款车】对比了昂克赛拉 起亚k3|朗动 轩逸 蓝鸟 朗逸这几款后 韩系车技术老旧被朋友给排除了；昂克赛拉虽然外观时尚 有创驰蓝天技术 但是自动挡要比卡罗拉贵2万 养护费用可能比卡罗拉要高 排除；轩逸和蓝鸟外配置相当 但新车没有啥优惠 排除；朗逸外观跟捷达一样 排除。最后在丰田故障率小 维护保养省钱 保值率高的口碑参考下选择了小卡。"|http://k.autohome.com.cn/spec/18890/view_1170228_1.html?st=112&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523175026|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 18:19:24|2016年06月26日 发表了口碑|来自：汽车之家iPhone版  2016年06月26日 发表了口碑  口碑   《卡罗拉的外观是我最看好的 当时再k3和卡罗拉做选选择》           【最满意的一点】手动档的车提速快 我喜欢提速的感觉 犀利的大灯 真是让人喜欢的不得了 我买的是外白内黑的 当时有一辆外白内黄的自动档的 我却没要【最不满意的一点】后来买完车交往了个女朋友 谁知媳妇的车是2011款马六 如果用两个车太浪费 她的怎么说也年岁久了 卖她那一部 可是我这个却是手动挡的 她说开着太费脑子 让现在的自动档气死了 以后大家谨记千万自动档 要不会有后悔的那天 开手动挡的 看着档次低【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】没有太中意的 直接看好这车了 直接去的莱州安利捷4s店【其他描述】|http://k.autohome.com.cn/spec/18891/view_1184866_1.html?st=10&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523176400|Autohome_review|뉴 보라(宝来)|ZHO|2016-06-27 18:19:26|2016年06月23日 发表了口碑|来自：手机汽车之家  2016年06月23日 发表了口碑  口碑   《稳固的德国工艺制作的底盘让弯道和颠簸路面不再那么困扰你。》   【最满意的一点】一般的油耗可以感受到大扭矩的动力。【最不满意的一点】内饰和外观设计中规中矩 想改装的部件较少。【空间】空间差异有点不足 宝来的价格桑塔纳的空间。【动力】动力杠杠的！宝来的价格近于高尔夫gti的享受【操控】前独立悬挂后连横式设计也是常规配置。【油耗】跟日系车没法比 相当于日系车安全性能也比不了一样。【舒适性】车内隔音效果相对比较不错的 【外观】个人比较喜欢外观改装的车型 宝来中规中矩外观改装的局限性很大。【内饰】座椅是高级仿pu的abs混合皮具 防龟裂较好 就是空间太不理想 宝来的价格桑塔纳的空间！【性价比】 总体来说宝来在同级车车里性价比很好 日系的卡罗拉ex 飞度 思域除了油耗低其他都是纸 韩系的k3 索纳塔 都是得个壳 国产的就不说了十几万买个国产仿制车没意思 法国和通用车那不是烧油是喝油。其他个各花入各眼【为什么最终选择这款车？】同价位的车对比中性价比很高 比国产 日 韩系车坚稳 比美国车省油。【其他描述】|http://k.autohome.com.cn/spec/14422/view_1181439_1.html?st=17&piap=0 633 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523200717|Autohome_review|랑동(朗动)|ZHO|2016-06-27 18:32:02|2016年06月21日 发表了口碑|来自：手机汽车之家  2016年06月21日 发表了口碑  口碑   《外观时尚好看 车子配置高实惠》           【最满意的一点】车子的外观和空间【最不满意的一点】1.6发动机动力不足【空间】后排虽然不能放倒 但足够日常生活所用 如何是放大东西的话就放不进去了【动力】起步肉 加速平稳 如果跑高速的话 油门响应有点慢 比如在跑高速过程中 你松下油门再想加速踩油门要踩深一点 中间有2秒的停顿加速【操控】方向盘轻 方向比较准【油耗】综合油耗还可以接受【舒适性】座椅很舒服 胎噪比较大跑高速【外观】外观非常喜欢【内饰】内饰中控台是软的比思域硬胶好很多【性价比】配置高 价格便宜实惠【为什么最终选择这款车？】选车中看了思域 速腾 卡罗拉 雷凌 k3。朗动的外观内饰价格优惠吸引我【其他描述】|http://k.autohome.com.cn/spec/20618/view_1178572_1.html?st=40&piap=0 2764 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523215541|Autohome_review|닛산 티아나(天籁)|ZHO|2016-06-27 18:41:01|2016年06月20日 发表了口碑|来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《性价比超高 外观大气稳重 省油。》             【最满意的一点】坐椅舒适 减震不错 空间宽敞 电动坐椅 后排出风口非常好。【最不满意的一点】自动大反应慢 基本没用 舒适版无倒车雷达 好歹十几万的车 居然不配这个两百块钱又非常实用的东西？前保险杠与叶子板接合处是水平状态 下雨天开车后污垢会从接合处流到保险杠上 很难看 我观察过其他车 其他车的这个部位一般都是有一个角度的 污水会顺着角度流到地上 不会弄脏保险杠 我认为这是设计不到位。【空间】很满意 现在看别人家的车都觉得小【动力】比原来的1.4强多了。【操控】没开过其他车 反正比k2好【油耗】没k2省 不过排量大0.6车重四百公斤 很不错了。我最低开过3.6升百公里 一般来说两百块跑四百三四十公里 高速城区农村各有一部分 如果纯城区只能跑三百六十左右。【舒适性】不错 买天籁就是冲这个来的 我腰椎间盘突出 做了手术 上了钢筋的 不能受冲击 过减速带比原来好多了【外观】大气稳重【内饰】还行 有味 但比原车好。【性价比】超高 别人都说这车得二十几万吧 我说十五万没人信。【为什么最终选择这款车？】由于前一个车是起亚k2 所以最先看的是k3 媳妇试坐之后认为除了大点之外和k2没啥区别 后来又试了一些其他车 都没感觉 直到走进一家店里看到天籁 媳妇坐进去试了一下 感觉很满意 移沙发确实不错 但是就是觉得价格超了 那是去年的事了 今年三月又去试了kx3 板车悬挂同样让人不满意 本地车展又去转了转 带媳妇去看了丰田卡罗拉 内饰丑死个人 比老款难看多了 后来媳妇发话 干脆一步到位 上天籁。【其他描述】|http://k.autohome.com.cn/spec/15104/view_1173431_1.html?st=54&piap=0 634 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523219452|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 18:43:01|2016年06月26日 发表了口碑|来自：汽车之家iPhone版  2016年06月26日 发表了口碑  口碑   《卡罗拉的外观是我最看好的 当时再k3和卡罗拉做选选择》           【最满意的一点】手动档的车提速快 我喜欢提速的感觉 犀利的大灯 真是让人喜欢的不得了 我买的是外白内黑的 当时有一辆外白内黄的自动档的 我却没要【最不满意的一点】后来买完车交往了个女朋友 谁知媳妇的车是2011款马六 如果用两个车太浪费 她的怎么说也年岁久了 卖她那一部 可是我这个却是手动挡的 她说开着太费脑子 让现在的自动档气死了 以后大家谨记千万自动档 要不会有后悔的那天 开手动挡的 看着档次低【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】没有太中意的 直接看好这车了 直接去的莱州安利捷4s店【其他描述】|http://k.autohome.com.cn/spec/18891/view_1184866_1.html?st=12&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523262177|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 19:09:01|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=165&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523262191|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 19:09:01|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=151&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523262215|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 19:09:01|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=129&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523262298|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 19:09:01|2016年06月19日 发表了口碑|来自：手机汽车之家  2016年06月19日 发表了口碑  口碑    《外观好看.性价比不错》             【最满意的一点】动力可以.颜值不错.空间杠杠的！油耗在接受范围内……不到五毛一公里.【最不满意的一点】避震较硬..隔音不太好..换档不是太顺..还有最重要的一点这款车居然只有一条智能钥匙.起亚有点抠哦！【空间】空间杠杠的.驾驶位我一米七的身高座的好宽松 特别是后座中间凸起几乎可以忽略 比帝豪强多了 帝豪后面凸起真心好高。【动力】对于在城里跑动力真心够用 如果不在乎油耗的话 只要舍得踩油门动力要多少是多少。【操控】指向没什么问题 就是方向盘有点重 换挡时有点卡 倒车时好容易熄火。六档位开起来好爽！【油耗】加了200跑了460多公里 算下来不到五毛一公里。油耗还是可以的 只是论坛里他们开出3～4毛一公里.所以觉得我的油耗还是下降空间滴！【舒适性】座椅还可以 就是隔音不是很好【外观】满分 开卡罗拉的朋友说我这张好有宽体轿跑的感觉??????【内饰】塑料感有点强【性价比】性价比没的说！非常可以！特别是15款！【为什么最终选择这款车？】最初是看上哈佛h5的 .奈何钱包米不够再加上我们当地的哈佛4s店服务真的太差了.直接是鼻子登天牛B哄哄的（昆明迪鑫）以后我还会买哈佛但绝对不在这家店买！不好意思情不自禁偏题了????言归正传 后来又去看远景看着看着就帝豪.看完后都决定上帝豪了.就在去订车的途中朋友说起他们店的15款k3在搞活动算下来跟帝豪差不多价格.然后就掉头直奔起亚家.直到定了车我才去论坛了解这款车.还好论坛里都说这张车不错【其他描述】把小三带回家绝不后悔 你值得拥有！导航和真皮座椅都是提车后在外面做的。|http://k.autohome.com.cn/spec/19723/view_1172428_1.html?st=67&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523262315|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 19:09:01|2016年06月20日 发表了口碑|来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《前脸16新款看上去比15款锐利了…》             【最满意的一点】最满意的就是性价比了…优惠过后同样的配置价格低…【最不满意的一点】提速有点慢…每次等红灯 都要深踩油门  中控丑 后备箱垫子塌陷…问4s怎么解决 竟然告诉我东西放两边 不要放中间 好吧 你赢了…【空间】对空间比较满意…媳妇说后排比她妹妹家索八小不多少…【动力】动力给4分吧 毕竟排量小…不过也够用了 【操控】没开过太多车 不懂操控 不过已经很满足了 操控比两轮电动车爽 哈哈…??【油耗】还在磨合期 上了高速匀速80 最低油耗5.2 比较满意吧【舒适性】前排舒适度不错…大儿子把后排当沙发蹦来蹦去…由此可见后面还是不错 【外观】这个要给满分 外表很漂亮 个人感觉比15款好看…【内饰】内饰只能给3分…虽然说看习惯了 但还是想说一句：太丑了…【性价比】性价比无敌…16增加了ESP 10.6万的车送了导航皮座椅贴膜脚垫…空间大 配置高 价格合适…总体来说还是瑕不掩瑜的…【为什么最终选择这款车？】选车历程比较艰辛…两个儿子了 用钱的地方太多 只有精打细算 虽然很想支持国产 但第一辆车还是打算耐用点 日系卡罗拉 1.6竟然没有ESP 而且价格偏高 美系新英朗 因为没买车之前用车都是借的表哥英朗 油耗有点高 也不想买同一个车了 别的就不说了 反正各种原因pass掉了 关注起亚其实是看中kx3了 无奈价格有点接受不了 前一段表妹家提了k3 感觉还不错 就把目光转投k3 事实证明车还是很不错的…【其他描述】喜欢就下手吧 普遍优惠都在1.5万左右 …不会让你失望的|http://k.autohome.com.cn/spec/25739/view_1174824_1.html?st=57&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523268272|Autohome_review|뉴 보라(宝来)|ZHO|2016-06-27 19:13:01|2016年06月23日 发表了口碑|来自：手机汽车之家  2016年06月23日 发表了口碑  口碑   《稳固的德国工艺制作的底盘让弯道和颠簸路面不再那么困扰你。》   【最满意的一点】一般的油耗可以感受到大扭矩的动力。【最不满意的一点】内饰和外观设计中规中矩 想改装的部件较少。【空间】空间差异有点不足 宝来的价格桑塔纳的空间。【动力】动力杠杠的！宝来的价格近于高尔夫gti的享受【操控】前独立悬挂后连横式设计也是常规配置。【油耗】跟日系车没法比 相当于日系车安全性能也比不了一样。【舒适性】车内隔音效果相对比较不错的 【外观】个人比较喜欢外观改装的车型 宝来中规中矩外观改装的局限性很大。【内饰】座椅是高级仿pu的abs混合皮具 防龟裂较好 就是空间太不理想 宝来的价格桑塔纳的空间！【性价比】 总体来说宝来在同级车车里性价比很好 日系的卡罗拉ex 飞度 思域除了油耗低其他都是纸 韩系的k3 索纳塔 都是得个壳 国产的就不说了十几万买个国产仿制车没意思 法国和通用车那不是烧油是喝油。其他个各花入各眼【为什么最终选择这款车？】同价位的车对比中性价比很高 比国产 日 韩系车坚稳 比美国车省油。【其他描述】|http://k.autohome.com.cn/spec/14422/view_1181439_1.html?st=18&piap=0 633 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523290095|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 19:28:01|2016年06月18日 发表了口碑|"2016年06月18日 发表了口碑  口碑    《空间大 省油 外观大气 优惠力度大》             【最满意的一点】空间大 油耗低 外观时尚 1万公里换机油保养。【最不满意的一点】没有ESP 没有发动机防盗 这俩项确实不应该简配。【空间】买车前参考过昂克赛拉 起亚k3|朗动 轩逸 蓝鸟 朗逸。轴距都是2700mm|但是看罗拉空间明显要大一些。180的大长腿坐进去都不挤。后排地面中间平整 也没有扶手 座三个175的壮汉也不觉得挤 不过后备箱不如轩逸的 感觉略小。【动力】1.6L的动力一个人开经常会有推背感 毕竟122马力 哈哈 但是座人了就感觉肉了 不过比朋友的斯柯达明锐1.6L双离合还是强劲不少 而且自然吸气的发动机跟涡轮增压比起来也没有烧机油的风险。【操控】之前开过面包车 开过荣威 但是跟卡罗拉的CVT比起来差远了 卡罗拉的标定确实比较扎实 换挡逻辑非常清新 开起来很平顺 出乎意料。在市区基本在1000转左右 处于ECO模式 高速跑120迈也就不到2000转左右 不知道需不需要像有的老司机说的过了磨合期高速拉缸。【油耗】刚提车时候油耗归零 开了110公里 竟然达到了惊人的4.1L/百公里 后来随着里程的增加逐步稳定在了6.5 6.6。日系车省油的名号确实不是盖的。【舒适性】这个价位的卡罗拉没有独立悬挂确实有些遗憾 在过减速带的时候 感觉略硬 风噪没有群友说的夸张 到了100迈内部还是比较安静的 但是偶尔能听到像石子刮地的声音 一直找不到原因。【外观】外观比老款的确实好看 个人觉得比雷凌的要收敛 离地间隙很低 好看但是也容易被磕碰。【内饰】内饰是硬塑料 黑白小仪表。10寸导航很加分 很大气 堪比K3.织物座椅去淘宝配个坐垫 美观舒适 朋友的真皮座椅夏天烫屁股。置物空间很多 放置杂物什么的没问题。【性价比】恰逢五一车展搞活动 优惠力度还是比较大了 送了贴膜导航装具行车记录仪。性价比相对来说要不算最好 中规中矩 总的来说推荐购买。【其它描述】没有ESP和自动落锁 后排座椅不能放倒......不能再多说了 毕竟才10万的合资车。【为什么最终选择这款车】对比了昂克赛拉 起亚k3|朗动 轩逸 蓝鸟 朗逸这几款后 韩系车技术老旧被朋友给排除了；昂克赛拉虽然外观时尚 有创驰蓝天技术 但是自动挡要比卡罗拉贵2万 养护费用可能比卡罗拉要高 排除；轩逸和蓝鸟外配置相当 但新车没有啥优惠 排除；朗逸外观跟捷达一样 排除。最后在丰田故障率小 维护保养省钱 保值率高的口碑参考下选择了小卡。"|http://k.autohome.com.cn/spec/18890/view_1170228_1.html?st=113&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523290384|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 19:28:01|2016年06月26日 发表了口碑|来自：汽车之家iPhone版  2016年06月26日 发表了口碑  口碑   《卡罗拉的外观是我最看好的 当时再k3和卡罗拉做选选择》           【最满意的一点】手动档的车提速快 我喜欢提速的感觉 犀利的大灯 真是让人喜欢的不得了 我买的是外白内黑的 当时有一辆外白内黄的自动档的 我却没要【最不满意的一点】后来买完车交往了个女朋友 谁知媳妇的车是2011款马六 如果用两个车太浪费 她的怎么说也年岁久了 卖她那一部 可是我这个却是手动挡的 她说开着太费脑子 让现在的自动档气死了 以后大家谨记千万自动档 要不会有后悔的那天 开手动挡的 看着档次低【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】没有太中意的 直接看好这车了 直接去的莱州安利捷4s店【其他描述】|http://k.autohome.com.cn/spec/18891/view_1184866_1.html?st=13&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523346888|Autohome_review|포커스(福克斯)|ZHO|2016-06-27 20:04:02|2016年06月20日 发表了口碑|"来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《唯一缺点就是空间小！》           【最满意的一点】好开 很稳 很省心 【最不满意的一点】空间小 降价快【空间】坐五个人不是太挤 后备箱比较大 综合还是不错【动力】不开空调 一个人开还是不错的 要舍得给油！驾驶乐趣不错 满座来空调那就力不从心了【操控】转向精准 悬架支撑不错 过弯比较有信心 过坑洼路面不是太舒服！【油耗】油耗还能接受 不是太高！当然没发和日系车比咯！【舒适性】座椅包裹性好 不过长途驾驶感觉不太舒服 座椅不是太软。关窗静音效果不错 胎噪有点大 其他方面都还不错的！【外观】外观还是比较漂亮的！轮毂再大一号就帅多了！【内饰】用料不错 做工就不敢恭维了！缝隙太大 不像合资的车。哎！真是应征了网友们所说的?百年福特毁于长安！希望长安福特之后们在做工方面改善改善！【性价比】性能不错 安全配置比较齐全 长安的价格贬值比较快！很让消费者伤心??买了车快两年了 唯一后悔的就是不该买最低配版的 如果再给我重新选择的机会 毫不犹豫直接上中高配！！！！！！！！！！【为什么最终选择这款车？】朗动 k3|朗逸。朗动挺漂亮 老婆看的时候说感觉太单薄.k3和朗动差不懂 配置也差不多 朋友的也是k3|不想大家都买一样的 果断放弃。朗逸神车 比较中庸 保值率高 不适合我们九零后 要有个性。福克斯基本安全配置比较高 油耗必上一代有所改善 车身扎实。比较适合自己 空间勉强够用 主要是自己开 能接受。【其他描述】油箱负压 空调效果不是很好 保养贵"|http://k.autohome.com.cn/spec/12132/view_1176643_1.html?st=112&piap=0 364 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523376176|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 20:23:03|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=167&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523376208|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 20:23:03|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=153&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523376626|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 20:24:09|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=131&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523376800|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 20:24:09|2016年06月19日 发表了口碑|来自：手机汽车之家  2016年06月19日 发表了口碑  口碑    《外观好看.性价比不错》             【最满意的一点】动力可以.颜值不错.空间杠杠的！油耗在接受范围内……不到五毛一公里.【最不满意的一点】避震较硬..隔音不太好..换档不是太顺..还有最重要的一点这款车居然只有一条智能钥匙.起亚有点抠哦！【空间】空间杠杠的.驾驶位我一米七的身高座的好宽松 特别是后座中间凸起几乎可以忽略 比帝豪强多了 帝豪后面凸起真心好高。【动力】对于在城里跑动力真心够用 如果不在乎油耗的话 只要舍得踩油门动力要多少是多少。【操控】指向没什么问题 就是方向盘有点重 换挡时有点卡 倒车时好容易熄火。六档位开起来好爽！【油耗】加了200跑了460多公里 算下来不到五毛一公里。油耗还是可以的 只是论坛里他们开出3～4毛一公里.所以觉得我的油耗还是下降空间滴！【舒适性】座椅还可以 就是隔音不是很好【外观】满分 开卡罗拉的朋友说我这张好有宽体轿跑的感觉??????【内饰】塑料感有点强【性价比】性价比没的说！非常可以！特别是15款！【为什么最终选择这款车？】最初是看上哈佛h5的 .奈何钱包米不够再加上我们当地的哈佛4s店服务真的太差了.直接是鼻子登天牛B哄哄的（昆明迪鑫）以后我还会买哈佛但绝对不在这家店买！不好意思情不自禁偏题了????言归正传 后来又去看远景看着看着就帝豪.看完后都决定上帝豪了.就在去订车的途中朋友说起他们店的15款k3在搞活动算下来跟帝豪差不多价格.然后就掉头直奔起亚家.直到定了车我才去论坛了解这款车.还好论坛里都说这张车不错【其他描述】把小三带回家绝不后悔 你值得拥有！导航和真皮座椅都是提车后在外面做的。|http://k.autohome.com.cn/spec/19723/view_1172428_1.html?st=69&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523376846|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 20:24:15|2016年06月20日 发表了口碑|来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《前脸16新款看上去比15款锐利了…》             【最满意的一点】最满意的就是性价比了…优惠过后同样的配置价格低…【最不满意的一点】提速有点慢…每次等红灯 都要深踩油门  中控丑 后备箱垫子塌陷…问4s怎么解决 竟然告诉我东西放两边 不要放中间 好吧 你赢了…【空间】对空间比较满意…媳妇说后排比她妹妹家索八小不多少…【动力】动力给4分吧 毕竟排量小…不过也够用了 【操控】没开过太多车 不懂操控 不过已经很满足了 操控比两轮电动车爽 哈哈…??【油耗】还在磨合期 上了高速匀速80 最低油耗5.2 比较满意吧【舒适性】前排舒适度不错…大儿子把后排当沙发蹦来蹦去…由此可见后面还是不错 【外观】这个要给满分 外表很漂亮 个人感觉比15款好看…【内饰】内饰只能给3分…虽然说看习惯了 但还是想说一句：太丑了…【性价比】性价比无敌…16增加了ESP 10.6万的车送了导航皮座椅贴膜脚垫…空间大 配置高 价格合适…总体来说还是瑕不掩瑜的…【为什么最终选择这款车？】选车历程比较艰辛…两个儿子了 用钱的地方太多 只有精打细算 虽然很想支持国产 但第一辆车还是打算耐用点 日系卡罗拉 1.6竟然没有ESP 而且价格偏高 美系新英朗 因为没买车之前用车都是借的表哥英朗 油耗有点高 也不想买同一个车了 别的就不说了 反正各种原因pass掉了 关注起亚其实是看中kx3了 无奈价格有点接受不了 前一段表妹家提了k3 感觉还不错 就把目光转投k3 事实证明车还是很不错的…【其他描述】喜欢就下手吧 普遍优惠都在1.5万左右 …不会让你失望的|http://k.autohome.com.cn/spec/25739/view_1174824_1.html?st=59&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
其他媒体|2523411214|bitauto|易车 > 问答 > 问题分类|ZHO|2016-06-27 20:45:02|东风悦达起亚k3码数拉不上怎么回事|东风悦达起亚k3码数拉不上怎么回事     提问者：易车网友 分类：  东风  其他  浏览[3]  2016-06-27 19:36  举报   东风悦达起亚k3码数拉不上怎么回事|http://ask.bitauto.com/detail/6709416/?leads_source=p029001|2016-06-27
기타|2523413720|Autohome_review|아반떼 AD(领动)|ZHO|2016-06-27 20:46:03|2016年06月02日 发表了口碑|来自：手机汽车之家  2016年06月02日 发表了口碑  口碑    《外观拉风 配置足够 整体性价比还是不错的。》           【最满意的一点】外观很拉风 现在路上还很少见 大轮毂。日间行车灯很高大上 自动头灯也很高端。中控台是软的 车内显示屏清晰度很高。倒车影像有随动辅助导线。很方便。车内音响很赞 我喜欢听音乐 完全满足我的要求。【最不满意的一点】后排不能放倒 这个真心很郁闷 这个放倒真的很难吗？这几天B柱内有异响 这还是新车呀 哎。。过几天去4s看看 希望不是啥大问题。另外胎噪确实大 我想跟轮胎大也有关系吧。悬挂还是有点硬 不过在接受范围内。【空间】空间同级别还是有优势的 中间无凸起。【动力】动力够用 现在用的eco模式【操控】转向精准 没啥虚位。【油耗】表显6 肯定是不准的 等下次油表亮再算算。【舒适性】还可以 家用够了。【外观】满意【内饰】做工还是比较好的 接缝均匀。【性价比】性价比高【为什么最终选择这款车？】同级别都看了 也试驾了 福克斯空间太小 科鲁兹都说油耗高 新英朗有点老气 卡罗拉没esp 思域根本没现车 看来看去家用也就韩系车了。【其他描述】换车的想法去年就有了 但是一直没有付诸行动 一是因为暂时有车开 二是今年上市新车多 想再等等 经常看论坛 心里已经有了几个备选 英朗 老表刚买的 开始觉得性价比很高 后来发现新旧差别很大 就pass了。福克斯外观不错 但是同事有好几辆 不想买一样的。k3性价比很高 优惠很大 但是新款感觉你没老款好看。看到最后就是领动了 配置高 外观拉风 总体性价比很高。|http://k.autohome.com.cn/spec/25701/view_1148059_1.html?st=115&piap=0 3959 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523413804|Autohome_review|아반떼 AD(领动)|ZHO|2016-06-27 20:46:04|2016年06月19日 发表了口碑|来自：手机汽车之家  2016年06月19日 发表了口碑  口碑    《选择不后悔 领动 领新而动。》             【最满意的一点】配置够用 外观造型动感。油耗表现好。磨合期过了后应该到正常水平了 现在降到8.3L了。【最不满意的一点】暂时还没发现 非要说的话速度上来后有点胎噪 另外轮胎有点卡小石子。【空间】我觉得空间很大了 后排的同事说不压抑 空间宽敞。头部空间和腿部空间都很充足 我身高173cm 不错。【动力】动力充足 只要肯给油 深踩油门 立马就走 反应灵敏 还没体验过运动模式 等磨合期完了试试。试驾的时候销售用1.4T的运动模式开过 感觉动力很猛。【操控】转向系统反应灵敏 方向盘虚位少 指向精准。悬架系统支撑性好 很稳。我在试驾的时候销售特地带我体验了一下转急弯 没有一点多余的倾斜。【油耗】刚提车的时候是18.几 慢慢的降下来了。满足预期 目前在磨合期 油耗下来了。【舒适性】座椅挺舒服的 我没加装真皮 感觉够用了。【外观】外观拉风 特别是前脸造型。【内饰】内饰设计很用心 能够平常接触的地方都是软材料 用心去体验啦。【性价比】自动精英版本配置够用了 具体的可以去看参数 选择不后悔。目前虽然没有大的降价 但是早买早享受了。【为什么最终选择这款车？】一直纠结着到底买哪款 去4s店看了好多车型 选车的时候看了卡罗拉 雷凌 起亚k3 领动 朗动 最终选择了领动 新款 1.6L购置税减半 自动精英型配置够用了。满意。另外就是感觉领动挺符合年轻人的气质的。我今年26岁 感觉其他车型不太符合 有的太中庸 有的太成熟了。这个刚刚好。还有就是胡歌代言的 挺喜欢胡歌的 哈哈 花痴了。【其他描述】今天看到了2辆白色的领动 对了 我定车那天4s店里的一台展车柠檬黄被人买了 很拉风。|http://k.autohome.com.cn/spec/25701/view_1171797_1.html?st=59&piap=0 3959 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523428442|Autohome_review|닛산 티아나(天籁)|ZHO|2016-06-27 20:55:02|2016年06月20日 发表了口碑|来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《性价比超高 外观大气稳重 省油。》             【最满意的一点】坐椅舒适 减震不错 空间宽敞 电动坐椅 后排出风口非常好。【最不满意的一点】自动大反应慢 基本没用 舒适版无倒车雷达 好歹十几万的车 居然不配这个两百块钱又非常实用的东西？前保险杠与叶子板接合处是水平状态 下雨天开车后污垢会从接合处流到保险杠上 很难看 我观察过其他车 其他车的这个部位一般都是有一个角度的 污水会顺着角度流到地上 不会弄脏保险杠 我认为这是设计不到位。【空间】很满意 现在看别人家的车都觉得小【动力】比原来的1.4强多了。【操控】没开过其他车 反正比k2好【油耗】没k2省 不过排量大0.6车重四百公斤 很不错了。我最低开过3.6升百公里 一般来说两百块跑四百三四十公里 高速城区农村各有一部分 如果纯城区只能跑三百六十左右。【舒适性】不错 买天籁就是冲这个来的 我腰椎间盘突出 做了手术 上了钢筋的 不能受冲击 过减速带比原来好多了【外观】大气稳重【内饰】还行 有味 但比原车好。【性价比】超高 别人都说这车得二十几万吧 我说十五万没人信。【为什么最终选择这款车？】由于前一个车是起亚k2 所以最先看的是k3 媳妇试坐之后认为除了大点之外和k2没啥区别 后来又试了一些其他车 都没感觉 直到走进一家店里看到天籁 媳妇坐进去试了一下 感觉很满意 移沙发确实不错 但是就是觉得价格超了 那是去年的事了 今年三月又去试了kx3 板车悬挂同样让人不满意 本地车展又去转了转 带媳妇去看了丰田卡罗拉 内饰丑死个人 比老款难看多了 后来媳妇发话 干脆一步到位 上天籁。【其他描述】|http://k.autohome.com.cn/spec/15104/view_1173431_1.html?st=55&piap=0 634 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523520980|Autohome_review|아반떼 AD(领动)|ZHO|2016-06-27 21:55:02|2016年06月02日 发表了口碑|来自：手机汽车之家  2016年06月02日 发表了口碑  口碑    《外观拉风 配置足够 整体性价比还是不错的。》           【最满意的一点】外观很拉风 现在路上还很少见 大轮毂。日间行车灯很高大上 自动头灯也很高端。中控台是软的 车内显示屏清晰度很高。倒车影像有随动辅助导线。很方便。车内音响很赞 我喜欢听音乐 完全满足我的要求。【最不满意的一点】后排不能放倒 这个真心很郁闷 这个放倒真的很难吗？这几天B柱内有异响 这还是新车呀 哎。。过几天去4s看看 希望不是啥大问题。另外胎噪确实大 我想跟轮胎大也有关系吧。悬挂还是有点硬 不过在接受范围内。【空间】空间同级别还是有优势的 中间无凸起。【动力】动力够用 现在用的eco模式【操控】转向精准 没啥虚位。【油耗】表显6 肯定是不准的 等下次油表亮再算算。【舒适性】还可以 家用够了。【外观】满意【内饰】做工还是比较好的 接缝均匀。【性价比】性价比高【为什么最终选择这款车？】同级别都看了 也试驾了 福克斯空间太小 科鲁兹都说油耗高 新英朗有点老气 卡罗拉没esp 思域根本没现车 看来看去家用也就韩系车了。【其他描述】换车的想法去年就有了 但是一直没有付诸行动 一是因为暂时有车开 二是今年上市新车多 想再等等 经常看论坛 心里已经有了几个备选 英朗 老表刚买的 开始觉得性价比很高 后来发现新旧差别很大 就pass了。福克斯外观不错 但是同事有好几辆 不想买一样的。k3性价比很高 优惠很大 但是新款感觉你没老款好看。看到最后就是领动了 配置高 外观拉风 总体性价比很高。|http://k.autohome.com.cn/spec/25701/view_1148059_1.html?st=118&piap=0 3959 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523521151|Autohome_review|아반떼 AD(领动)|ZHO|2016-06-27 21:55:02|2016年06月19日 发表了口碑|来自：手机汽车之家  2016年06月19日 发表了口碑  口碑    《选择不后悔 领动 领新而动。》             【最满意的一点】配置够用 外观造型动感。油耗表现好。磨合期过了后应该到正常水平了 现在降到8.3L了。【最不满意的一点】暂时还没发现 非要说的话速度上来后有点胎噪 另外轮胎有点卡小石子。【空间】我觉得空间很大了 后排的同事说不压抑 空间宽敞。头部空间和腿部空间都很充足 我身高173cm 不错。【动力】动力充足 只要肯给油 深踩油门 立马就走 反应灵敏 还没体验过运动模式 等磨合期完了试试。试驾的时候销售用1.4T的运动模式开过 感觉动力很猛。【操控】转向系统反应灵敏 方向盘虚位少 指向精准。悬架系统支撑性好 很稳。我在试驾的时候销售特地带我体验了一下转急弯 没有一点多余的倾斜。【油耗】刚提车的时候是18.几 慢慢的降下来了。满足预期 目前在磨合期 油耗下来了。【舒适性】座椅挺舒服的 我没加装真皮 感觉够用了。【外观】外观拉风 特别是前脸造型。【内饰】内饰设计很用心 能够平常接触的地方都是软材料 用心去体验啦。【性价比】自动精英版本配置够用了 具体的可以去看参数 选择不后悔。目前虽然没有大的降价 但是早买早享受了。【为什么最终选择这款车？】一直纠结着到底买哪款 去4s店看了好多车型 选车的时候看了卡罗拉 雷凌 起亚k3 领动 朗动 最终选择了领动 新款 1.6L购置税减半 自动精英型配置够用了。满意。另外就是感觉领动挺符合年轻人的气质的。我今年26岁 感觉其他车型不太符合 有的太中庸 有的太成熟了。这个刚刚好。还有就是胡歌代言的 挺喜欢胡歌的 哈哈 花痴了。【其他描述】今天看到了2辆白色的领动 对了 我定车那天4s店里的一台展车柠檬黄被人买了 很拉风。|http://k.autohome.com.cn/spec/25701/view_1171797_1.html?st=62&piap=0 3959 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523600912|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 22:46:01|2015年10月15日 发表了质量评价|2015年10月15日 发表了质量评价  质量   【车身外观】  侧滑门-门把手或门锁(扣)操控困难  【行驶过程】  刹车时(车身)会振动-在低速刹车时        2015年08月08日 发表了口碑  口碑    《两年前就心有所属 喜欢k3 不后悔》             【最满意的一点】乘坐空间和舒适性都还不错 外观和内饰设计在同级别也都还好【最不满意的一点】暂时还没有发现【空间】比较好 后排前排都不错【动力】觉得挺好 超车也快【操控】中规中矩 家用车【油耗】目前还没有降下去 在使用一段时间【舒适性】挺好 坐过的人都说好【外观】看个人喜好 我很喜欢【内饰】整体做工还不错 中控像驾驶员侧倾斜 不错【性价比】整体不错【其它描述】人无完人 车无完车 我觉得车也是有生命的 要好好待它【为什么最终选择这款车】喜欢3有两年了 一见钟情 现在终于实现了  第一次看见3儿[色] 是2013年的时候 当时没想那么多就是觉得好看 当时我的大学生涯才开始一半 不管是在家的这座城市还是上学的那座城市 走在街上遇到3儿都会多看两眼 慢慢的 两年多已经过去了 3儿虽不是什么豪车 但是我感觉就像一个亲人一样 脑子里只要是关于车的方面 3儿就会第一时间浮现 从未改变过[微笑]。 上学的时候只是心里偶尔想过[害羞] 如果我将来经济独立了 肯定会买这个车 未必买好车 但是要买合适的 当时同学嘴里说的都是豪车[撇嘴] 我只是淡淡一笑 觉得他们的梦想是好的 但是我更喜欢切合实际[微笑]。 到了今年2015年 终于毕业了[害羞] 回到了家里的城市 运气好 工作也算稳定。每天基本也会是家--单位。[糗大了] 家里有个06年12月出产的伊兰特 每次洗干净 感觉也挺好 主要我也爱收拾 别人都说这车最多两年吧 ^_^ 有些得意[得意] 现在毕业工作了 我爸爸和我单位又没在一起 哎 这下可咋办[可怜]你们懂得[坏笑]开过的车也不少 B50、景程、雅阁、智跑、高尔夫、2000、捷达、福克斯、速腾、CRV、翼虎、k2、赛欧等等。虽然都不是些豪车[嘘] 但咱也只是平常老百姓呀[委屈] [嘘]告诉你们个秘密 现在经常去健身房 因为3儿很美 我就是为了和3儿 以后看起来更和谐 不能胖开着它呀[害羞] 7月最后一个星期 打算去离我们最近的一个4S店哄背ぞ眉⒖闯担20多公里路程吧 没想到去了以后顺带订车。[阴险][阴险][阴险]最后的结果是手动GLS 送皮座椅 氙灯 侧厚膜 挡泥板..101000 唉就这样了 勉强能接受 最后落地114000多 希望大家有时间都来临潼玩儿 这里有什么 你们自己去百度 不会让你们失望滴我还算是个对生活有规划的人 15年前半年目前有了3儿 工作也还算稳定 家庭比较和谐美满。希望后半年会有一个女朋友 和我相遇、相知、相爱、相伴、相守 然后走进婚姻的殿堂。希望也会有喜欢这个车的女孩 一定也非常美...[害羞] 等有了女朋友后 想再发一个媳妇儿当车模 到时候兄弟们多多鼓励支持呀[抱拳][抱拳]|http://k.autohome.com.cn/spec/19723/view_700200_1.html?st=168&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523600939|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 22:46:01|2016年06月04日 发表了口碑|来自：手机汽车之家  2016年06月04日 发表了口碑  口碑   《外观漂亮 内饰不错 油耗可以接收 胎噪有点大》           【最满意的一点】外观漂亮 感觉比朗动耐看 内饰看着舒服【最不满意的一点】胎噪很大 很烦人 没esp.esp.esp.重要事情说三遍 为啥国内生产的车不能标配 也用不了多少成本 【空间】够大 家用没问题【动力】一般【操控】还能接受【油耗】一般【舒适性】较硬【外观】漂亮【内饰】漂亮 做工也可以【性价比】挺高【为什么最终选择这款车？】看了 本田凌派 现代朗动 丰田卡罗拉 雷凌 开始最钟意本田凌派 1.8排量没有购置税减半政策 所以放弃 现代朗动外形漂亮 接受不了内饰 放弃 不喜欢卡罗拉外形 中网像个小胡子 和雷凌一样 内饰看着不像10万的车 放弃 无意间看见k3 外形够漂亮 内饰好看 韩国车这几年进步还是挺快的【其他描述】|http://k.autohome.com.cn/spec/25737/view_1149586_1.html?st=154&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523600993|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 22:46:01|2016年06月08日 发表了追加口碑|2016年06月08日 发表了追加口碑 追加    购车1年7个月后追加口碑    当前行驶里程 17500 公里 当前平均油耗 7.0 升/百公里    免费保养 1 次  收费保养 4 次  共花费 526.00 元   【油耗】东风悦达起亚k3的油耗总体来说还行不耗油 但也不是特别省油对1.6排量的车来说只能是说的过去 1年6个月综合油耗7.0到7.5之间 但感觉不是很准确有偏差。【保养】保养多是按保养手册全部4s店5000公里保养一次 价格还可以接受 到目前为止只做常规保养 我选用了道达尔的机油发动机声音小加速有力跟同级别比【故障】故障率到目前为止就两个 一个启动机得问题冷车启动异响批次问题已经解决 还一个就是车身异响问题 特别是b柱一到冬天的时候就响 应该是热胀冷缩的 也还可以接受不打算拆 怕拆了后有后遗症。【吐槽】当然也是要吐槽一下的 也10多万的车了音响主机能不能换好点 跟面包车一样一点多没有听歌乐趣 说是有6个喇叭 但跟4个喇叭没有什么区别那个音质 还有那个车内气味太大了不好散掉 多快2年的车了味道还是很大时间久了头痛 不会甲醛超标吧 还一个减震问题 开起来没有舒适感 还没有面包车舒服就是一个硬 还有一个灯光问题太差了实在是太差了 虽然近光带透镜但亮光也太差了吧 在城市里面还能勉强一上高速就危险了 害的还要自己在掏钱换灯泡无语了 但k3这个我买的不后悔 它的优点多过缺点 从来没有把我丢在路上之少但目前来说是这样 之后会怎么样只能走一步算一步|http://k.autohome.com.cn/spec/19724/view_581942_1.html?st=132&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523601138|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 22:46:01|2016年06月19日 发表了口碑|来自：手机汽车之家  2016年06月19日 发表了口碑  口碑    《外观好看.性价比不错》             【最满意的一点】动力可以.颜值不错.空间杠杠的！油耗在接受范围内……不到五毛一公里.【最不满意的一点】避震较硬..隔音不太好..换档不是太顺..还有最重要的一点这款车居然只有一条智能钥匙.起亚有点抠哦！【空间】空间杠杠的.驾驶位我一米七的身高座的好宽松 特别是后座中间凸起几乎可以忽略 比帝豪强多了 帝豪后面凸起真心好高。【动力】对于在城里跑动力真心够用 如果不在乎油耗的话 只要舍得踩油门动力要多少是多少。【操控】指向没什么问题 就是方向盘有点重 换挡时有点卡 倒车时好容易熄火。六档位开起来好爽！【油耗】加了200跑了460多公里 算下来不到五毛一公里。油耗还是可以的 只是论坛里他们开出3～4毛一公里.所以觉得我的油耗还是下降空间滴！【舒适性】座椅还可以 就是隔音不是很好【外观】满分 开卡罗拉的朋友说我这张好有宽体轿跑的感觉??????【内饰】塑料感有点强【性价比】性价比没的说！非常可以！特别是15款！【为什么最终选择这款车？】最初是看上哈佛h5的 .奈何钱包米不够再加上我们当地的哈佛4s店服务真的太差了.直接是鼻子登天牛B哄哄的（昆明迪鑫）以后我还会买哈佛但绝对不在这家店买！不好意思情不自禁偏题了????言归正传 后来又去看远景看着看着就帝豪.看完后都决定上帝豪了.就在去订车的途中朋友说起他们店的15款k3在搞活动算下来跟帝豪差不多价格.然后就掉头直奔起亚家.直到定了车我才去论坛了解这款车.还好论坛里都说这张车不错【其他描述】把小三带回家绝不后悔 你值得拥有！导航和真皮座椅都是提车后在外面做的。|http://k.autohome.com.cn/spec/19723/view_1172428_1.html?st=70&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523601156|Autohome_review|K3(起亚K3)|ZHO|2016-06-27 22:46:01|2016年06月20日 发表了口碑|来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《前脸16新款看上去比15款锐利了…》             【最满意的一点】最满意的就是性价比了…优惠过后同样的配置价格低…【最不满意的一点】提速有点慢…每次等红灯 都要深踩油门  中控丑 后备箱垫子塌陷…问4s怎么解决 竟然告诉我东西放两边 不要放中间 好吧 你赢了…【空间】对空间比较满意…媳妇说后排比她妹妹家索八小不多少…【动力】动力给4分吧 毕竟排量小…不过也够用了 【操控】没开过太多车 不懂操控 不过已经很满足了 操控比两轮电动车爽 哈哈…??【油耗】还在磨合期 上了高速匀速80 最低油耗5.2 比较满意吧【舒适性】前排舒适度不错…大儿子把后排当沙发蹦来蹦去…由此可见后面还是不错 【外观】这个要给满分 外表很漂亮 个人感觉比15款好看…【内饰】内饰只能给3分…虽然说看习惯了 但还是想说一句：太丑了…【性价比】性价比无敌…16增加了ESP 10.6万的车送了导航皮座椅贴膜脚垫…空间大 配置高 价格合适…总体来说还是瑕不掩瑜的…【为什么最终选择这款车？】选车历程比较艰辛…两个儿子了 用钱的地方太多 只有精打细算 虽然很想支持国产 但第一辆车还是打算耐用点 日系卡罗拉 1.6竟然没有ESP 而且价格偏高 美系新英朗 因为没买车之前用车都是借的表哥英朗 油耗有点高 也不想买同一个车了 别的就不说了 反正各种原因pass掉了 关注起亚其实是看中kx3了 无奈价格有点接受不了 前一段表妹家提了k3 感觉还不错 就把目光转投k3 事实证明车还是很不错的…【其他描述】喜欢就下手吧 普遍优惠都在1.5万左右 …不会让你失望的|http://k.autohome.com.cn/spec/25739/view_1174824_1.html?st=60&piap=0 2886 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523608888|Autohome_review|뉴 보라(宝来)|ZHO|2016-06-27 22:50:06|2016年06月23日 发表了口碑|来自：手机汽车之家  2016年06月23日 发表了口碑  口碑   《稳固的德国工艺制作的底盘让弯道和颠簸路面不再那么困扰你。》   【最满意的一点】一般的油耗可以感受到大扭矩的动力。【最不满意的一点】内饰和外观设计中规中矩 想改装的部件较少。【空间】空间差异有点不足 宝来的价格桑塔纳的空间。【动力】动力杠杠的！宝来的价格近于高尔夫gti的享受【操控】前独立悬挂后连横式设计也是常规配置。【油耗】跟日系车没法比 相当于日系车安全性能也比不了一样。【舒适性】车内隔音效果相对比较不错的 【外观】个人比较喜欢外观改装的车型 宝来中规中矩外观改装的局限性很大。【内饰】座椅是高级仿pu的abs混合皮具 防龟裂较好 就是空间太不理想 宝来的价格桑塔纳的空间！【性价比】 总体来说宝来在同级车车里性价比很好 日系的卡罗拉ex 飞度 思域除了油耗低其他都是纸 韩系的k3 索纳塔 都是得个壳 国产的就不说了十几万买个国产仿制车没意思 法国和通用车那不是烧油是喝油。其他个各花入各眼【为什么最终选择这款车？】同价位的车对比中性价比很高 比国产 日 韩系车坚稳 比美国车省油。【其他描述】|http://k.autohome.com.cn/spec/14422/view_1181439_1.html?st=19&piap=0 633 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523622826|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 22:59:01|2016年06月18日 发表了口碑|"2016年06月18日 发表了口碑  口碑    《空间大 省油 外观大气 优惠力度大》             【最满意的一点】空间大 油耗低 外观时尚 1万公里换机油保养。【最不满意的一点】没有ESP 没有发动机防盗 这俩项确实不应该简配。【空间】买车前参考过昂克赛拉 起亚k3|朗动 轩逸 蓝鸟 朗逸。轴距都是2700mm|但是看罗拉空间明显要大一些。180的大长腿坐进去都不挤。后排地面中间平整 也没有扶手 座三个175的壮汉也不觉得挤 不过后备箱不如轩逸的 感觉略小。【动力】1.6L的动力一个人开经常会有推背感 毕竟122马力 哈哈 但是座人了就感觉肉了 不过比朋友的斯柯达明锐1.6L双离合还是强劲不少 而且自然吸气的发动机跟涡轮增压比起来也没有烧机油的风险。【操控】之前开过面包车 开过荣威 但是跟卡罗拉的CVT比起来差远了 卡罗拉的标定确实比较扎实 换挡逻辑非常清新 开起来很平顺 出乎意料。在市区基本在1000转左右 处于ECO模式 高速跑120迈也就不到2000转左右 不知道需不需要像有的老司机说的过了磨合期高速拉缸。【油耗】刚提车时候油耗归零 开了110公里 竟然达到了惊人的4.1L/百公里 后来随着里程的增加逐步稳定在了6.5 6.6。日系车省油的名号确实不是盖的。【舒适性】这个价位的卡罗拉没有独立悬挂确实有些遗憾 在过减速带的时候 感觉略硬 风噪没有群友说的夸张 到了100迈内部还是比较安静的 但是偶尔能听到像石子刮地的声音 一直找不到原因。【外观】外观比老款的确实好看 个人觉得比雷凌的要收敛 离地间隙很低 好看但是也容易被磕碰。【内饰】内饰是硬塑料 黑白小仪表。10寸导航很加分 很大气 堪比K3.织物座椅去淘宝配个坐垫 美观舒适 朋友的真皮座椅夏天烫屁股。置物空间很多 放置杂物什么的没问题。【性价比】恰逢五一车展搞活动 优惠力度还是比较大了 送了贴膜导航装具行车记录仪。性价比相对来说要不算最好 中规中矩 总的来说推荐购买。【其它描述】没有ESP和自动落锁 后排座椅不能放倒......不能再多说了 毕竟才10万的合资车。【为什么最终选择这款车】对比了昂克赛拉 起亚k3|朗动 轩逸 蓝鸟 朗逸这几款后 韩系车技术老旧被朋友给排除了；昂克赛拉虽然外观时尚 有创驰蓝天技术 但是自动挡要比卡罗拉贵2万 养护费用可能比卡罗拉要高 排除；轩逸和蓝鸟外配置相当 但新车没有啥优惠 排除；朗逸外观跟捷达一样 排除。最后在丰田故障率小 维护保养省钱 保值率高的口碑参考下选择了小卡。"|http://k.autohome.com.cn/spec/18890/view_1170228_1.html?st=114&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523623099|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-06-27 22:59:01|2016年06月26日 发表了口碑|来自：汽车之家iPhone版  2016年06月26日 发表了口碑  口碑   《卡罗拉的外观是我最看好的 当时再k3和卡罗拉做选选择》           【最满意的一点】手动档的车提速快 我喜欢提速的感觉 犀利的大灯 真是让人喜欢的不得了 我买的是外白内黑的 当时有一辆外白内黄的自动档的 我却没要【最不满意的一点】后来买完车交往了个女朋友 谁知媳妇的车是2011款马六 如果用两个车太浪费 她的怎么说也年岁久了 卖她那一部 可是我这个却是手动挡的 她说开着太费脑子 让现在的自动档气死了 以后大家谨记千万自动档 要不会有后悔的那天 开手动挡的 看着档次低【空间】【动力】【操控】【油耗】【舒适性】【外观】【内饰】【性价比】【为什么最终选择这款车？】没有太中意的 直接看好这车了 直接去的莱州安利捷4s店【其他描述】|http://k.autohome.com.cn/spec/18891/view_1184866_1.html?st=14&piap=0 526 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523637025|Autohome_review|랑동(朗动)|ZHO|2016-06-27 23:07:49|2016年06月21日 发表了口碑|来自：手机汽车之家  2016年06月21日 发表了口碑  口碑   《外观时尚好看 车子配置高实惠》           【最满意的一点】车子的外观和空间【最不满意的一点】1.6发动机动力不足【空间】后排虽然不能放倒 但足够日常生活所用 如何是放大东西的话就放不进去了【动力】起步肉 加速平稳 如果跑高速的话 油门响应有点慢 比如在跑高速过程中 你松下油门再想加速踩油门要踩深一点 中间有2秒的停顿加速【操控】方向盘轻 方向比较准【油耗】综合油耗还可以接受【舒适性】座椅很舒服 胎噪比较大跑高速【外观】外观非常喜欢【内饰】内饰中控台是软的比思域硬胶好很多【性价比】配置高 价格便宜实惠【为什么最终选择这款车？】选车中看了思域 速腾 卡罗拉 雷凌 k3。朗动的外观内饰价格优惠吸引我【其他描述】|http://k.autohome.com.cn/spec/20618/view_1178572_1.html?st=41&piap=0 2764 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523683884|Autohome_review|랑동(朗动)|ZHO|2016-06-27 23:38:02|2016年06月21日 发表了口碑|来自：手机汽车之家  2016年06月21日 发表了口碑  口碑   《外观时尚好看 车子配置高实惠》           【最满意的一点】车子的外观和空间【最不满意的一点】1.6发动机动力不足【空间】后排虽然不能放倒 但足够日常生活所用 如何是放大东西的话就放不进去了【动力】起步肉 加速平稳 如果跑高速的话 油门响应有点慢 比如在跑高速过程中 你松下油门再想加速踩油门要踩深一点 中间有2秒的停顿加速【操控】方向盘轻 方向比较准【油耗】综合油耗还可以接受【舒适性】座椅很舒服 胎噪比较大跑高速【外观】外观非常喜欢【内饰】内饰中控台是软的比思域硬胶好很多【性价比】配置高 价格便宜实惠【为什么最终选择这款车？】选车中看了思域 速腾 卡罗拉 雷凌 k3。朗动的外观内饰价格优惠吸引我【其他描述】|http://k.autohome.com.cn/spec/20618/view_1178572_1.html?st=42&piap=0 2764 0 0 2 0 0 0 0 0 1|2016-06-27
기타|2523690802|Autohome_review|포커스(福克斯)|ZHO|2016-06-27 23:43:02|2016年06月20日 发表了口碑|"来自：手机汽车之家  2016年06月20日 发表了口碑  口碑    《唯一缺点就是空间小！》           【最满意的一点】好开 很稳 很省心 【最不满意的一点】空间小 降价快【空间】坐五个人不是太挤 后备箱比较大 综合还是不错【动力】不开空调 一个人开还是不错的 要舍得给油！驾驶乐趣不错 满座来空调那就力不从心了【操控】转向精准 悬架支撑不错 过弯比较有信心 过坑洼路面不是太舒服！【油耗】油耗还能接受 不是太高！当然没发和日系车比咯！【舒适性】座椅包裹性好 不过长途驾驶感觉不太舒服 座椅不是太软。关窗静音效果不错 胎噪有点大 其他方面都还不错的！【外观】外观还是比较漂亮的！轮毂再大一号就帅多了！【内饰】用料不错 做工就不敢恭维了！缝隙太大 不像合资的车。哎！真是应征了网友们所说的?百年福特毁于长安！希望长安福特之后们在做工方面改善改善！【性价比】性能不错 安全配置比较齐全 长安的价格贬值比较快！很让消费者伤心??买了车快两年了 唯一后悔的就是不该买最低配版的 如果再给我重新选择的机会 毫不犹豫直接上中高配！！！！！！！！！！【为什么最终选择这款车？】朗动 k3|朗逸。朗动挺漂亮 老婆看的时候说感觉太单薄.k3和朗动差不懂 配置也差不多 朋友的也是k3|不想大家都买一样的 果断放弃。朗逸神车 比较中庸 保值率高 不适合我们九零后 要有个性。福克斯基本安全配置比较高 油耗必上一代有所改善 车身扎实。比较适合自己 空间勉强够用 主要是自己开 能接受。【其他描述】油箱负压 空调效果不是很好 保养贵"|http://k.autohome.com.cn/spec/12132/view_1176643_1.html?st=113&piap=0 364 0 0 2 0 0 0 0 0 1|2016-06-27
其他媒体|1644663996|mobile01|新進文章|ZHO|2015-02-05 00:12:01|關於HD PENTAX-DA 16-85mm....|"本來小弟打算自己打一篇文不過上網找資料時發現這位前輩文筆甚好早已回答了小弟心中的疑問又提出更多精闢見解在徵得對方同意之後(感謝Waltyu兄無私分享）於此登出全文及其鏈結小弟僅將Waltyu兄的分析加上紅色以利閱讀無更改任何內容（有的話請告知小弟改正）希望可以提供眾壇友另一個面相來討論這顆新鏡頭原文聯結以下為原文Mobile 01「防塵防滴搭載 兼顧輕量與小廣角‧HD PENTAX-DA 16-85mm F3.5-5.6 ED DC WR」全破解以文找文waltyu 在天空部落發表於17:12:47   Pentax專欄 作為第一篇中文的Pentax DA16-85的測試 m01網站的測試報告引起了Pentax使用者的不少迴響。但打從民國89年當時打著「華人最大」的攝影家手札就發生過對大眾品牌和小眾品牌的測試報告立場不公的情形。於是先有Minolta Fan Club後有Pentax Fan Club的誕生。現在臉書上一些創作者很容易遭到不同政治立場的網軍檢舉 維護自己言論自由的基本方是就是「向臉書買廣告」當保險 這樣就不會動不動被檢舉到下架。同樣地 如果Pentax總代理富堃也有這種敏銳度 相信m01的測試報告就不會在Pentax設群中引起軒然大波。以下為本人就該篇測試報告的破解http://www.mobile01.com/newsdetail.php?id=16222原文「Ricoh在Photokina 2014一共展示了三顆新鏡頭 而這三顆鏡頭當中也只有HD PENTAX-DA 16-85mm F3.5-5.6 ED DC WR公佈正式的鏡頭規格 其它兩顆鏡頭分別會是恆定光圈的中望遠變焦鏡以及高望遠變焦鏡頭 至於詳細規格還是得等到原廠宣布。HD PENTAX-DA 16-85mm F3.5-5.6 ED DC WR的出現其實很難去界定它在K接環所扮演的角色的角色 因為上有smc PENTAX-DA 18-135mm F3.5-5.6 ED AL[IF] DC WR下有smc PENTAX-DA 17-70mm F4AL[IF] SDM 兩者分別具備7.5x光學變焦以及f/4恆定光圈的優勢 所以我想HD PENTAX-DA 16-85mm F3.5-5.6 ED DC WR只是提供消費者更多元的選擇 等效24mm的廣角端、新加入的HD 多層鍍膜、WR耐候能力 在未來可能會作為Kit鏡也說不定。」 分析1：DA16-85的定位非常明確 就是入門級變焦(DA18-55)、中階變焦(DA17-70)、高階變焦(DA★16-50|DA20-40LE)和高倍率變焦鏡(DA18-135|DA18-270)中的中階變焦鏡頭。中階鏡頭畫質比入門級鏡頭和旅遊鏡佳 方便性比高階鏡頭佳（廣角更廣 望遠更遠） 其定位非常明確。DA16-85很明顯是取代DA17-70的 除非DA17-70也改款為HD DA17-70WR 否則「只是提供消費者更多元的選擇」這個論點是缺乏基本觀念下自己硬套的解釋！DA17-70在DA16-85推出後說穿了已經沒有市場 個人認為在庫存清倉完後官網就會移入停產商品類別 也就是說生產線實際已經停產 只是還有庫存。 「新中階標準變焦鏡」的定位在明顯不過！ 你會說Canon在EF-S17-85IS之後推出EF-S15-85IS是「只是提供消費者更多元的選擇」嗎？EF-S15-85當然是EF-S17-85的後繼款阿 DA16-85和DA17-70的關係也一樣 m01這位編輯的水準光第一段就表露無遺了。原文 「上圖是HD PENTAX-DA 16-85mm F3.5-5.6 ED DC WR鏡頭的正面及背面 鏡身外觀雖然是塑膠材質 但整體處理的還不錯亦不會有廉價感 反而這顆鏡頭的價格讓人有點摸不著頭緒 日本官網上的價格￥80|600（含稅） 怎麼算都超過新台幣兩萬元 以鏡頭規格與用料來看 這價格並不怎麼友善 預計會比富堃官網上的DA 18-135mm F3.5-5.6及DA17-70mm F4貴上至少7000元！但新鏡總是有蜜月期的 不急的話倒是可以等價格趨近穩定 或是其它用戶的評價再做打算。」 分析2：我們來比較一下Canon|Nikon同級鏡的價格 以日本原廠建議售價為準 因為Canon官網只有未稅價 故均以未稅價比較。Pentax DA16-85WR ￥74|630 Nikon AF-S16-85VR ￥95|000Canon EF-S15-85IS ￥105|000加上固定比例的消費稅(也就是我國的營業稅)後價格高低順序並不會因此改變。 注意這三款鏡頭中Nikon是最早發表的 另外Canon也已經過了剛發售價格最高的時期(這裡是指市場實際售價 與前面的官方建議售價無關)。但是新上市Nikon可以賣貴 Canon可以賣貴 Pentax卻不能賣貴 這樣論述公平嗎？(剛上市價格高對廠商來講也是利用想搶鮮的客戶願意多負一點錢來加速回收研發成本) 用料的部分Pentax 12群16枚（非球面鏡片3枚、ED鏡片1枚）Nikon 11群17枚（非球面鏡片3枚、ED鏡片2枚）Canon 12群17枚（非球面鏡片3枚、UD鏡片1枚）有明顯不如C|N嗎？原文「這顆鏡頭在前玉部分有加上SP鍍膜 目的就是提供更防油防水的保護能力 但這鍍膜可不是無敵...因為再怎麼厲害還是無法防刮 另外鍍膜也是有壽命的 長時間擦拭鍍膜還是會被消耗殆盡 建議還是乖乖買一片保護鏡比較實在。」分析3：這段很有趣………Pentax官網http://www.ricoh-imaging.co.jp/japan/products/lens/technology/SP（Super Protect）コーティングSPコーティング撥水性、撥油性にすぐれたペンタックス独自の特殊コーティング。高性能レンズの第１面に採用し、レンズ面の保護に効果を発揮しています。このコーティングはホコリや水滴、油などがつきにくいだけでなく、万一汚れが付着した場合にも、簡単に落としやすいという特長をそなえています。Pentax官網沒有介紹影片 但可以參考下列實測影片https://www.youtube.com/watch?v=ZIlUwfhKAwA Nikon官網http://www.nikon-image.com/products/lens/about/technology.htmlフッ素コート【Fluorine Coat】汚れが付着しにくく付着しても簡単に拭き取れるニコンのフッ素コートは、優れた防汚性能でレンズ表面に汚れ（埃、水滴、油、泥）が付着しにくく、付着した場合も簡単に拭き取り可能です。しかも、ニコン独自のコーティングテクノロジーで、耐久性が極めて高くコーティングが剥がれにくいため、他の同様のコーティングよりもはるかに多くの拭き取り回数に耐え、その優れた効果が長期にわたって持続します。反射防止効果もあり、クリアーな画像の撮影にも貢献します。AF-S NIKKOR 400mm f/2.8E FL ED VR、AF-S NIKKOR 300mm f/4E PF ED VR、AF-S TELECONVERTER TC-14E IIIに採用しています。Canon官網http://cweb.canon.jp/ef/technology/eflens-technology.htmlフッ素コーティングフッ素コーティングレンズ表面に付着した汚れを簡単に取り除くことを目的として開発された新しいコーティング技術。それが、フッ素コーティングです。撥油性・撥水性が高く、溶剤を使わずに乾いた布で取り除くことが可能。乾拭き後に静電気を帯びにくく、ホコリなどを寄せ付けにくいのも特長です。表面が滑らかで傷つきにくく、水滴がつきにくい特性もあります。 Nikon和Canon稱為氟鍍膜 Pentax則沒有說明SP鍍膜的成分 不過其實都是抗污防潑水鍍膜。Pentax是第一個推出的 因此除了第一批發表的少數幾款DA鏡頭(例如DA14|DA40LE|DA16-45)之外幾乎都有SP鍍膜。Canon和Nikon都是近年才推出的(Pentax現在官網能查到最早的鏡頭是97年 但實際上更早) Canon只有L鏡才有 像EF24F2.8IS|EF35F2.0IS這種鏡頭都沒有 Pentax則是DA35F2.4|DA50F1.8都有。Nikon則是只有三款鏡頭有 Nikon的宣傳影片看起來可能效果更勝SP鍍膜 但SP鍍膜一來是推出時間早 二來是普及率高 可以得知Pentax和Canon|Nikon的想法不同 C|N要多花點錢買高階鏡頭才能享受到抗污防潑水鍍膜 Pentax則是很容易就享受到。 M01有本事的話等AF-S NIKKOR 300mm f/4E PF ED VR的測試文也來寫「這顆鏡頭在前玉部分有加上SP鍍膜 目的就是提供更防油防水的保護能力 但這鍍膜可不是無敵...因為再怎麼厲害還是無法防刮 另外鍍膜也是有壽命的 長時間擦拭鍍膜還是會被消耗殆盡 建議還是乖乖買一片保護鏡比較實在。」這種廢話給大家瞧瞧 說m01沒有品牌本位主義嗎？你相信？ 原文「HD PENTAX-DA 16-85mm F3.5-5.6 ED DC WR的焦段涵蓋廣角與中望遠 等效焦長為24.5-130mm 換算下來約5.3倍光學變焦 美中不足的當然還是那個光圈大小 如果是f/2.8起跳或許會更有吸引力。鏡片結構採12群16枚的設計 其中包括了三枚非球面鏡片以及一枚ED超低色散鏡片 另外「HD鍍膜」的加入更是這顆鏡頭的重點 而HD鍍膜也就是SMC的進化版 而這些搭載HD鍍膜的新鏡頭在外觀最不一樣的地方就是捨棄過去的SMC的「綠圈」塗裝 用「紅圈」作為HD鍍膜的識別方式 且日後也不再會有SMC新鏡的出現 因為原廠已經確定停產了 這是2013年就公佈的訊息 相信一些老用戶淚都已經流乾了吧。至於HD鍍膜所強調的優勢就是在逆光環境下可以盡可能避免眩光、鬼影的產生 雖然SMC鍍膜在過去就是以抗耀光的能力著稱 或許HD鍍膜的表現更上層樓 另外對畫質也有提升 特別是提升影像的銳利度與對比度 另外就是散景比過去的SMC鍍膜柔和 不過最後這點則是見仁見智 畢竟每個人看散景的標準不盡相同。此外目前的HD鏡頭都改用圓形光圈 過去的多邊形光圈設計恐怕要成為歷史。」分析3：嫌最大光圈沒有F2.8 難道Canon|Nikon有16-85F2.8了嗎？Sigma|Tamron|Tokina至今也沒有這種產品。在底片時代只有Minolta AF24-105F3.5-4.5是望遠端超過85mm且最大光圈維持F4.5 像Nikon AF-D24-120F3.5-5.6和Tamron SP24-135F3.5-5.6望遠端光圈都是F5.6 這種情況至今沒有打破 拿一款沒有一個品牌有出的規格來嫌Pentax 憑空想想真是好棒棒！ 再來 第一款HD鏡頭是101年9月11日發表的HD DA560http://www.ricoh-imaging.co.jp/japan/news/2012/********_7.html「同一天」也發表了smc DA18-270http://www.ricoh-imaging.co.jp/japan/news/2012/********_9.html 此外 上個月才在CES展上展示搭配K-50後繼機的新入門級標準變焦鏡 就是smc DA L18-50F4-5.6https://www.flickr.com/photos/scott_burnham/***********/http://news.ricoh-imaging.co.jp/rim_info/2015/********_006329.html信口開河寫測試文真是不負責任！原文 「這張也是用最短對焦距離35公分拍攝的成果 很可惜放大倍率不夠 不然這樣的焦段又能兼具微距功能的話 吸引力肯定會更大。」分析4：最高放大倍率與最近對焦距離Pentax最近對焦距離35cm最高放大倍率0.26XNikon最近對焦距離38cm最高放大倍率1/4.6(0.217X)Canon最近對焦距離35cm最高放大倍率0.21X M01是在拐灣罵AF-S16-85VR和EF-S15-85IS放大倍率不夠嗎？Pentax可是三款鏡頭中最高放大倍率最高的喔！原文 「DA在Pentax代表的是數位專用鏡 所以在鏡身上看不到光圈環的結構 不過很可惜的是連對焦視窗或是對焦距離的符號提示都沒有 以兩萬多元的鏡頭來說 這樣的設計還挺沒有誠意的。」分析5：沒有對焦距離視窗的批評是正確的 但是什麼年代了還在講光圈環？原文 「雖然K3推出至今已有一年多的時間 但它目前還是Pentax在數位單眼相機領域的機皇 當然還是選擇它來搭配HD PENTAX-DA 16-85mm F3.5-5.6 ED DC WR 而且K3的耐候能力在業界也有極高的評價。其實小編自己也猜不透為什麼Penatx遲遲不推出全片幅數位單眼相機 旗下有一堆鏡頭根本就是為全片幅量打造 但用戶卻苦無解放的機身 直到最近我才晃然大悟 因為Penatx把眼光放得更遠 直接挑戰中片幅相機 就像是去年推出的645Z 其感光元件尺寸是35mm全片幅的1.7倍 畫質在國內外都獲得許多專業攝影師的推崇 重點是它的價格才23萬出頭 在以C/P來說在中片幅領域幾乎找不到對手 同時還有機會吸引到35mm全片幅的用戶 因為單純就畫素跟畫質來看的話 645Z應該是完勝目前的35mm機種 日後若有機會也會進行645Z的測試 敬請期待！」分析6：1.現有的FA鏡頭只有FA31LE|FA43LE|FA77LE|FA35|FA50 DFA鏡頭只有DFA50macro|DFA100macro 要推35mm數位單眼非常缺鏡頭是原廠多年來數次在訪談中清楚說明的事實。2.看起來這位編輯居然連Pentax在底片時代就有做645相機都不知道。 原文「以上是鏡頭廣角端與望遠端鏡頭伸出後的差異 這顆鏡頭採外變焦內對焦的結構 也就是說變焦時鏡頭長度會變化 而對焦時鏡頭長度不會改變亦不會旋轉 如此一來搭配偏光鏡作業時就不會受到影響；此外HD PENTAX-DA 16-85mm F3.5-5.6 ED DC WR支援全時手動對焦 在半按快門合焦成功後 維持半按快門的動作同時可以調整對焦環來選擇你所需要的對焦距離。以下緊接著就是一連串的光學品質測試 對這顆新鏡頭有興趣的朋友可別錯過了。」分析7:Pentax的Quick-shift focus system不是真正的全時手動對焦 這位編輯的中文程度需要加強。原文 「這顆新鏡在畫質上的表現有點讓我訝異 簡單來說廣角端中央畫質從開放光圈就很銳利 不過邊緣畫質從開放光圈到最小光圈都屬於不及格狀態。中央畫質從f/3.5到f/11的表現都很好 而從上圖妳可以發現f/16開始出現衰退情形 當光圈縮到最小f/22時候畫質也顯得最差；但是邊緣畫質從f3.5開始就糊的非常誇張 就算是f/8的表現也只稱得上堪用 小編原本還懷疑是不是指定的裁切區域有問題 但把原圖放大到100%仔細端詳一番才知道 測試過程本身以及裁切區域並沒有問題 而是影像中央以外1/2的畫質的確是有待改善。」分析8：這大概可以說是網路上的測試的通病。鏡頭在設計時檢查中央和邊緣畫質 用的測試圖表是平面的還是立體的大家可以想想看 有的鏡頭像場平整 有的鏡頭全開的景深是一個弧形 既然是用這種非「固定測試場景」的測試 確實是可以反應實際拍攝遇到的情形 但是難道如果換C|N的測試 場景又變了 這種結果可以拿來比較嗎？P|N|C都有公布MTF 如果P被講成這麼差 用同樣的標準那C|N又會好到哪去？ Pentax DA16-85http://www.ricoh-imaging.co.jp/japan/products/lens/k/standard/hdpentax-da-16-85/Nikon AF-S16-85http://www.nikon-image.com/products/lens/nikkor/af-s_dx_nikkor_16-85mm_f35-56g_ed_vr/spec.htmlCanon EF-S15-85http://cweb.canon.jp/ef/lineup/ef-s/ef-s15-85-f35-56/spec.html原文 「望遠端的表現可就好多了 讓我們從中央畫質開始看起 從f/5.6到f/11之間的畫質都還不錯 f/16可以發現畫質有了輕微的變化 f/22開始出現衰退的情形直到最小光圈 而f/40的中央畫質我個人則是完全無法接受 看起來就像是未合焦的影像；邊緣畫質f/8到f/16是我唯一可以接受的範圍 其餘之外的畫質都是鬆散到不行。」分析9：筆者拍照超過15年 從來沒用過F40拍照 如果讀者有這種癖好 K-3在v1.10版韌體中也首創「繞射補償」 今天換AF-S16-85或EF-S15-85 不要說同樣F40畫質有差多少 C|N的機身可以做數位繞射補償？顯然這位編輯完全不知道K-3有這項獨步武林的功能。http://www.ricoh-imaging.co.jp/japan/support/download/digital/k3_s.html 原文「16mm廣角端拍攝：這顆鏡頭內含三枚非球面鏡片 而非球面鏡片的目的就是改善像差及變形 但從實際拍攝的結果來看 表現似乎是差強人意 等效24.5mm的桶狀變形非常明顯 但這是為經機身數位修正後的表現 因為K3韌體目前還不支援 只能等日後更新再看看修正的幅度了。」分析10：如果Pentax的標準稱為「差強人意」 那Sony Vario-Sonnar T*16-80F3.5-4.5ZA這款還掛卡爾蔡司的叫？http://www.photozone.de/sony-alpha-aps-c-lens-tests/141-zeiss-za-16-80mm-f35-45-dt--sony-alpha--review--test-report?start=1原文 「自從HD鍍膜加入後 這類鏡頭的另一個特性就是採用圓形光圈 意指縮光圈之後拍攝得到的散景也會是圓形 這顆鏡頭的光圈由七枚光圈葉片組成 以星芒公式來看可獲得14道星芒角 而有趣的是從開放光圈就可以看到星芒角的出現但有點偏細 f/5.6-f/8的星芒則是有點發育不良的感覺 f/11你會發現星芒角會有分叉的情況 最討喜的時刻我想就是在f/22的時候 因為看起來比較健康」分析11：真是隨便寫隨便錯 DA★55F1.4SDM就是smc鍍膜但有圓形光圈的。圓形光圈的定義是指「從最大光圈到縮1.5-2（依品牌及款式不同）級後散景維持圓形」。還有底片時代沒有人在講星芒 底片時代有需要的話有星芒鏡（濾鏡）。原文 「這款新鏡頭最特別的地方就是加入HD鍍膜 而HD鍍膜以官方的定義來說 目的就是擁有更出色的抗耀光能力 盡可能的抑制眩光及鬼影 但從實測結果來看好像不是這麼回是...從f/5.6就出現了明顯的光斑 縮1又1/3級光圈光斑就誇張成這樣...光圈繼續縮下去的表現想必更慘 我想各位從上圖的測試結果已經可以得到答案 以上是擷取照片中央1/2的影像 需要檢視原圖的話建議下載壓縮檔。」分析12：抗耀光一向是Pentax在日系品牌中 「要是Pentax說自己是第二 沒有人敢講自己是第一」的情況 m01既然把Pentax講成這麼爛 那就拿C|N也在同樣情況下PK一下看看鹿死誰手阿。原文 「約一週左右的時間試用下來 我必須很誠實的告訴各位 這顆鏡頭的C/P值並不高 且大部分的表現都只能說是中規中矩 雖然偶有佳作出現但也的確只是小小的亮點 並不會讓你有衝動敗家的慾望 而這個亮點就是散色的抑制能力 另外就是無須特別縮光圈在中央畫質就能有不錯的表現 但前提是你必須忍受影像邊緣那鬆散卻又無可救藥的畫質 其實從原廠的MTF來看應該沒那麼誇張 但實際測出來的結果卻是如此 這讓小編感到有些懊惱 因為這是我第一次遇到在縮光圈之後邊緣畫質還不見提升的鏡頭 但尷尬的就是它又稱得上是一顆旅遊鏡 風景題材的拍攝也絕對少不了 但要風景攝影玩家接受中央以外的影像畫質不佳可能不是一件容易的事情 畢竟這不是大光圈鏡頭 就算邊緣畫質不好我也可以善用大光圈優勢讓影像邊緣畫質不佳的部分給柔化掉。 改紅圈之後的HD鍍膜沒有想像中厲害是我意料之外的事情 因為這不就是它主打的特色嗎？怎麼一測就崩壞了...對焦速度是我個人滿在意的部分 就算搭配K3這類高階機種 其實對焦速度也不算快 當然這是小編使用過眾多品牌、機型後所得到的結論 畢竟它也稱不上高階鏡頭 這樣的表現我並不意外。24.5-130mm的等效焦長在構圖取景時還算是方便 比較可惜的就是放大倍率不夠 只有0.26x而已連拍小花或桌上的美食都有吃力。這顆鏡頭在小編眼中雖然差強人意 不過這或許是各位期待已久的焦段或是規格 畢竟K-Mount可用的副廠鏡頭實在有限 用戶們不是彼此交流二手鏡 就是只能存錢等待貴鬆鬆的新鏡頭 若你對HD PENTAX-DA 16-85mm F3.5-5.6 ED DC WR還有期待的話 不妨參考文末更多的實拍範例 謝謝各位。」分析13:結論 看了這麼多跟本是浪費生命阿！這種帶有品牌成見的文章如果不是要寫破解我還真沒興趣花時間去看。DA20-40LE一年前剛上市時價格也是比較高 但現在水貨的價格只要兩萬初就有了 那個品牌不是剛上市很貴一年後會降價？一款鏡頭以撰稿者的水準用一週就能徹底體會體會它的品質？筆者一直不談邊角畫質的問題 最主要是因為筆者沒沒無名不像m01隨便就可以跟代理商借到鏡頭。DA18-135的邊角畫質就真的是不太理想（但不是全焦段 各種距離都有這種情況） 看了前面那麼多偏頗的論述 對邊角畫質這點……看看日本Map Camera的測試…….國內流水帳的測試隨便看看就算了吧。http://news.mapcamera.com/KASYAPA.php?itemid=26117&catid=281"|http://www.mobile01.com/topicdetail.php?f=251&t=4260364|2015-02-05
各大媒体|1644941855|gmw|滚动读报|ZHO|2015-02-05 05:41:02|k3s最高降1.7万元|"*************-02-05 04:32:42.0k3s最高降1.7万元k3s;最高;降;1.7;万;元********滚动读报/enpproperty-->url:http://epaper.jinghua.cn/html/2015-02/05/content_170440.htm|id:0京华时报讯（记者麦田）上周六 记者从东风悦达起亚经销商处了解到 起亚k3s最高可享1.5万元现金优惠 置换购车还可享受5000元置换补贴。据经销商介绍 由于k3s上市以来一直保持了不错的销量 此前很长一段时间k3s的优惠幅度徘徊在1.2万元上下 近期价格继续下探 最高降价幅度达到1.5万元。据了解 k3s需求量较大的车型为1.6升gl自动挡 指导价11.18万元 降价幅度为1.4万元 优惠后售价为9.78万元；指导价14.38万元的1.6升premium自动挡车型可优惠1.7万元 优惠后售价12.68万元。据悉 k3s共有6款车型在售 均搭载1.6升排量的发动机。目前自动挡车型现车相对较多 颜色以黑、白为主 但1.6升两款手动挡车型现车很少 个别颜色需要预订 定金2000元 两周左右可提车。"|http://news.gmw.cn/newspaper/2015-02/05/content_104338042.htm|2015-02-05
各大媒体|1676796776|12365auto|质量投诉|ZHO|2015-02-26 10:30:02|2015款东风悦达起亚K3冷启动异响|投诉编号：【84123】 投诉品牌： 东风悦达起亚 投诉车系： 起亚K3 投诉车型： 2015款 1.6L 手动 GLS 投诉时间： 2015-2-25 22:30:14    投诉内容： 天气冷的时候冷启动时发动机舱传出“扑哧“的一声 很刺耳 自己录的音和视频4s店不认可 要他们自己听到才诊断 但是那声音时有时无 去4s店100多公里。已经有很多k3车主遇到了这个问题 都是起动机复位不及时造成的 并已经更换起动机 为什么厂家就没有别的方法诊断呢？非要听到那异响声才肯更换起动机呢？本来就是车子质量问题还没有一个比较简单的处理方式 这样就变相增加了车主开支(过路费 油费 住宿费)。那厂家除了更换起动机其他费用就该车主自己承担吗？   投诉回复： 中国汽车质量网已将您的投诉转给生产企业以及政府有关主管部门 我们将会对此投诉继续跟踪 请您持续关注！|http://www.12365auto.com/zlts/20150225/84123.shtml|2015-02-26
其他媒体|1676956373|zhidao_baidu|生活|ZHO|2015-02-26 12:06:02|比亚迪k3怎么关收音机||http://zhidao.baidu.com/question/1755458631770165988.html?entry=qb_browse_default|2015-02-26
汽车社区|1677394451|autohome_cn|狮跑论坛|ZHO|2015-02-26 16:49:01|起亚 皮卡 很酷！有没有？（附KIA历史）|2011-8-9 11:51:49    起亚 皮卡 很酷！有没有？（附KIA历史）        简介        起亚汽车（Kia Motors）是现代起亚汽车集团的子公司 也是韩国第二大汽车制造商 总部位于首尔。起亚汽车是韩国最老牌的汽车公司。1944年底 二战还没有结束 势衰力竭的日军还没有完全撤离朝鲜半岛。在12月的一天 起亚公司的前身京城精工终于突破种种困难在汉城成立了 对于每个起亚人甚至整个韩国汽车工业来说 这一时刻是值得纪念的。 历程  起亚成立于1944年 是韩国历史最悠久的汽车公司 原本是由制造钢管和自行车起家。1952年 起亚开始生产摩托车、卡车和房车。七、八十年代 起亚受惠于亚洲经济起飞 规模不断扩大 并于1986年开始冲出海外。1992年起亚进军美国市场 短短数年在美国各地已都有其代理商出售起亚汽车。然而 亚洲金融风暴爆发波及韩国 起亚在1997年破产 导致起亚51%股权被转手到其国内对手──现代汽车。后来现代公司重组 目前现代汽车公司已拥有起亚40%股权。当时 韩国国内的经济和工业百废待兴 多年的战火洗礼使韩国人民生活水平已经接近了最低标准 汽车在当时还是件奢侈的玩意。当年京城精工所生产的是流行的代步工具--脚踏车。1945年初 生产脚踏车的工厂已初具规模 到第二年春天 韩国国内第一款脚踏车出厂。之后的15年中 公司一直默默生产他们的脚踏车 同时投入利润不断扩大工厂规模。1960年工会成立后不久 公司决定生产他们的第一种摩托化产品 而被命名c-100的摩托车在1961年10月正式出厂 第二年 一辆小型的厢式三轮货车k360也面世。从此 起亚走上了“automobile”之路。1971年 起亚服务公司成立 开始对已经大量售出的三轮货车提供保障 并且有意发展四轮汽车 毕竟这是公司发展和壮大的必然路径。同年公司推出四轮厢式货车titan。由于当时韩国经济的飞速发展 这种轻型的多用途货车非常受一些刚开始创业的小公司和个体户青睐 销量急速攀升。1974年 公司第一辆采用汽油发动机的小型轿车brisa诞生 从此 起亚开始与世界车厂的发展方向接轨 并且介入竞争激烈的轿车市场之中。1975年 brisa的皮卡版本b-1000出厂 没多久 起亚就推出了一款新车--k303 这款家庭轿车与十分稚嫩的brisa相比有明显的进步和成熟 所以取得较大的销售效益。但是 由于多种原因 起亚当时生产的轿车还存在明显的缺陷 加上在新车型的开发设计上出现了问题 公司决定首先要借鉴国外行进车型生产的成功经验。于是在1979年 起亚仿制了法国标志 的604轿车 并且组装了意大利菲亚特的132型轿车。        为了公司的长远发展 1984年 起亚r&d中心正式建立 肩负起起亚汽车的技术研究和新产品开发设计的任务 为日后起亚公司丰富完善的车型体系和先进的科技含量打下坚实基础 同时也坚定了起亚“走自己路”的决心。1986年 起亚自行设计的小型乘用车brisa出厂 同年起亚与美国福特汽车公司达成合作协议 并且开始设计和生产采用了福特技术的pride车型。1988年 rhino和trade两款厢式货车出厂 标志着公司在大力发展轿车的同时仍然对货车生产给予高度重视。1989年7月 起亚在东京建立了研究院 4个月后 起亚经济研究中心也宣告成立。进入九十年代 起亚有了一项很大的改变。1990年3月 公司正式改名为起亚汽车株式会社(kia motors corporation) 紧接着亚山湾工厂竣工 之后 potentia、sephia和sportage等车型陆续出现 起亚进入了发展的黄金时期。1994年 起亚公司度过了自己的50岁金禧盛典 但公司的经营出现了问题 发展令人担忧。在国内和北美这两个起亚的最大市场上 销售成绩不断下滑 起亚r&d中心也由于资金问题不得不关闭。1996年 起亚公司作出了购买英国莲花公司小型开蓬跑车elan生产权的决定 并且由起亚自行对该车作出修改 以适应相对的客户群。可惜这辆漂亮的小车却胎死腹中 没生产几辆就被搁置了。  另：东风悦达起亚汽车有限公司系由东风汽车公司、江苏悦达投资股份有限公司、韩国起亚自动车株式会社共同组建的中外合资轿车制造企业。 所属子品牌 ： 霸锐 Borrego (大型SUV)欧菲莱斯 Opirus佳乐 Carens索兰托 Sorento (中大型SUV)欧迪玛 Optima (中型家庭房车)帝国 Imperial首都 Capital狮跑 Sportage (小型SUV)克利多斯 Credos普莱特 Pride锐欧 Rio (小型五人车)    [ 本帖最后由 foryou97 于 2011-08-09 11:57:18 编辑 ]     用户名   操作   操作时间   查看全部|http://club.autohome.com.cn/bbs/thread-c-565-11661571-1.html|2015-02-26
其他媒体|1778118614|hexun|滚动新闻 > 全部新闻|ZHO|2015-04-30 18:32:01|起亚k3s到底怎么样 悦达起亚k3s报价 起亚k3s口碑 起亚k3s全国最低价|"　　北京博润中信汽车销售有限公司东风悦达起亚4s店发布：起亚K3S现车齐全 继续底价促销 综合优惠可达4万元。购车可享受免费新车检测 代办临牌 汽车交强险商业险等业务 另外还可免费获赠原厂DVD导航 全车贴膜 封釉封塑 发动机护板 地胶 大包围脚垫 麂皮 掸子 香水 把套等万元精美汽车装饰礼包。此活动面对全国 感兴趣的各地新老客户可垂询热线：*********** 曹经理 （全国销售热线）　　车型名称厂商指导价现价优惠幅度现车情况2014款起亚K3S 1.6L 手动GL10.18万6.184万有现车2014款起亚K3S 1.6L 自动GL11.18万7.184万有现车2014款起亚K3S 1.6L 手动GLS11.48万7.484万有现车2014款起亚K3S 1.6L 自动GLS12.48万8.484万有现车2014款起亚K3S 1.6L 自动DLX13.18万9.184万有现车2014款起亚K3S 1.6L 自动Premium14.38万10|384万有现车　　K3S独有的运动风格、高标准的安全性和尖端的科技配备 为您打造独一无二的尊贵气质。动感激情、活力四射的肆意驰骋 与您的风格品味相得益彰。狭长的虎啸式前中网承袭起亚家族特征 张扬的进气格栅 打造出令人过目不忘的“吞噬感” 更显时尚运动。K3S丰富多彩的空间性 多样式座椅折叠功能 超强货物容纳能力 保障安全、便利的驾驶。K3S安装了以性能为中心的高效技术的发动机让驾驶者在无论何种路况能感受运动风格的驾驶体验 尽享驰骋的快感。　　北京博润中信汽车销售有限公司-东风悦达起亚 4S 店提供了很多附加增值性服务 如直赔保险和贷款 下表将为您提供更多有用信息：起亚K3S车型在该店的保养、贷款、保险情况保养信息质保期5年或100000公里店内建议保养周期7500公里更换机油机滤费用600元左右　　(以4S店价格为准)更换机油三滤费用800元左右　　(以4S店价格为准)保险信息店内提供保险公司人保保险费用5500元左右　　(以4S店价格为准)　　编辑点评：　　K3S是东风悦达起亚最新推出的一款紧凑运动型车。该车全系只搭载1.6L自然吸气发动机 最大功率128马力 峰值扭矩156牛・米 匹配6速手自一体变速箱或6速手动变速箱。经销商名称：北京博润中信汽车销售有限公司联系电话:*********** 曹经理公司地址：北京市北五环仰山桥往北天通苑 （地铁5号线天通苑站)　　如系本站原创文章 转载请注明出处：汽车中国。（责任编辑：HN666）"|http://auto.hexun.com/2015-04-30/175456752.html|2015-04-30
其他媒体|1778267619|hexun|滚动新闻 > 全部新闻|ZHO|2015-04-30 20:13:01|2015款起亚k3多少钱 无底线优惠价格 销售全国 全新优惠 报价及图片|　　北京博润中信汽车销售有限公司东风悦达起亚4s店发布：起亚K3现车充足 继续底价促销 综合优惠可达4万元。购车可享受免费新车检测 代办临牌 汽车交强险商业险等业务 另外还可免费获赠原厂DVD导航 全车贴膜 封釉封塑 发动机护板 地胶 大包围脚垫 麂皮 掸子 香水 把套等万元精美汽车装饰礼包。此活动面对全国 感兴趣的各地新老客户可垂询热线：*********** 曹经理 （全国销售热线）　　起亚K3 相关配置及报价车型指导价(万)4s店价格(万)价格变化(万)备注1.6L 手动GL10.286.28↓4现车1.6L 自动GL11.287.28↓4现车1.6L 手动GLS11.487.48↓4现车1.6L 自动GLS12.488.48↓4现车1.6L 自动DLX13.189.18↓4现车1.6L 自动Premium14.3810.38↓4现车1.8L 自动Premium14.9814.58↓4现车全国销售热线：*********** 曹经理　　k3在前脸的设计上十分突出力量感和线条的精炼 采用起亚旗舰车型K9的镀铬直瀑式竖条进气格栅 视觉感受更为大气、稳健 后尾组合尾灯和外后视镜集成转向灯都采用LED设计 再配合LED日间行车灯 彰显出浓厚的科技感以及时代感 在精炼线条勾勒下 大倾角前风挡以及溜背式车尾处理都传递出独特的动态肌肉造型美 视觉冲击强烈 很容易给人留下深刻的印象。　　K3还搭载了起亚最新的1.6L伽马D-CVVT和1.8L Nu D-CVVT两款发动机 最大功率分别达到128马力和146马力 动力强劲且燃油经济性突出。配合先进的6速手自一体变速箱 操控随心 能很好的开发车主驾驭热情。安全方面 K3很好的继承了K系家族优良的安全传统 以C-NCAP全新五星标准打造 搭配了VSM车辆动态控制系统、6方位安全气囊 TPMS胎压监测、HID氙气大灯、前后泊车辅助系统等高科技配置。起亚K3在4S店部分保养信息保养消息质保周期5年或者10万公里店内建议保养周期3个月或者5000公里更换机油机滤费用322元更换机油三滤费用汽滤价格=机油两滤价格+150左右　　注：以上部分价格会与实际情况有差异 真实价格以到店为准。制表：汽车中国　　起亚K3以新颖的外形和丰富的配置引来不少消费者的关注。起亚K3不但在舒适性配置上更加丰富 而且主动安全性也得到了提升。目前 店内起亚K3现车销售 购车最高优惠4万元 店内还提供了各种金融贷款方案。感兴趣的朋友可到店或电话咨询。经销商名称：北京博润中信汽车销售有限公司联系电话:***********曹经理公司地址：北京市北五环仰山桥往北天通苑 （地铁5号线天通苑站)　　如系本站原创文章 转载请注明出处：汽车中国。（责任编辑：HN666）|http://auto.hexun.com/2015-04-30/175459657.html|2015-04-30
其他媒体|1799598393|zhidao_baidu|生活|ZHO|2015-05-14 08:29:01|朗动科鲁兹雷凌k3优缺电点|来自：手机知道互联网|http://zhidao.baidu.com/question/682390672245092812.html?entry=qb_browse_default|2015-05-14
其他媒体|1825426770|hexun|滚动新闻 > 全部新闻|ZHO|2015-05-29 10:04:01|15款奥迪A3现车最高优惠8万全国上牌|　　奥迪A3 准确的说是一汽-大众奥迪A3 2014年上市以来一直都以符合国人审美观念的外观、简约而又不简单的内饰以及出色的动力表现深受消费者的青睐。近日 小编从北京博奥众诚汽车销售有限公司　　了解到 15款奥迪A3月底冲量 现车最高优惠8万元 可全国上牌 手续齐全 感兴趣的朋友可以致电经销商以便了解更多详情。　　具体车型售价见下表：车型厂家指导价经销商报价优惠幅度Limousine40TFSI自动豪华型29.67万21.67万80000元Sportback35TFSI手动进取型18.49万11.49万70000元Sportback35TFSI自动进取型19.99万12.99万70000元　　制表：汽车中国 http://carschina.com注：车辆价格随时变化 敬请随时关注当地市场　　外观方面 奥迪A3与A4L的设计中饱含了一辆运动型轿车惯有的组合元素。高挑的侧面腰线巧妙连接着头尾灯组 使车身整体感更加强烈 结合了外扩的轮拱造型 动感气质油然而生 镀铬边框装点下的侧窗形态使得这两款车型在视觉效果上显得分外协调。　　内饰方面 全新A3采用了非常简洁的内饰设计 位于中控台顶部是一款可升降的7英寸液晶显示屏 可显示行车电脑、蓝牙电话及音响系统。中控台控制面板仅存几个功能按键 让日常操作变得简单 中控台顶部由大面积的软性材质覆盖 手感还算不错。　　编辑点评：　　全新国产奥迪A3与现款相比在尺寸上已经进行了超越 三门版达到了2601mm、五门版为2650mm。但即便如此 五门版奥迪A3相比奔驰全新B级、宝马全新1系也依然处于劣势地位。喜欢这款车的朋友可以来电（店）了解咨询。　　注文章内的价格为编辑在“市场前线”真实采集到的当日价格 由于汽车价格变化多端 同时此价格是经销商的个体行为 所以价格仅供参考使用。另外 文中图片为车型资料片 价格信息与图片拍摄地点无关。　　更多详情请联系经销商：公司名称:北京博奥众诚汽车销售有限公司经营性质: 综合联系人:张先生销售电话:***********E-mail:**********@qq.com公司网址:http://www.im4s.cn/30981地址:北京市朝阳区立水桥北苑路93号报上您是来自于“汽车中国网站”的用户 将会得到更多的优惠　　如系本站原创文章 转载请注明出处：汽车中国。（责任编辑：HN666）|http://auto.hexun.com/2015-05-29/176286898.html|2015-05-29
其他媒体|1826037198|hexun|滚动新闻 > 全部新闻|ZHO|2015-05-29 16:37:04|北京起亚K3全系最高优惠5万 销售全国 起亚K3最新报价表 优惠详情 性能评测|"　　起亚k3最高优惠4万元 并有全车2万精品装饰赠送 目前店内有现车充足 颜色齐全 对该车感兴趣的朋友可致电经销商详询。24小时热线电话：*********** 张经理　　起亚K3最新报价表车型(北京报价)指导价(万)4s店价格(万)价格变化(万)备注1.6L 手动GL2014款10.287.283现车1.6L 自动GL2014款11.288.283现车1.6L 手动GLS2014款11.488.484现车1.6L 自动GLS2014款12.489.484现车1.6L 自动DLX2014款13.1810.184现车1.6L 自动Premium2014款14.3811.384现车1.8L 自动Premium2014款14.9811.984现车24小时热线电话：*********** 张经理　　K3是起亚家族中全新的一款紧凑型家轿 一经推出就以其前卫时尚的外形 在年轻消费群体中拥有了较高人气。车型配置丰富 空间实用 油耗适中 适合一般家庭使用。不足之处：动力不足 底盘偏软 操控性一般 定价偏高。　　北京地区 东风悦达起亚4S店提供了很多附加增值性服务 如直赔保险和贷款 下表将为您提供更多有用信息请您参考：起亚K3车型在该店的保养、贷款、保险情况保养信息质保周期三年或10万公里店内建议保养周期5000公里更换机油机滤费用　　350元左右　　（以4S店价格为准）更换机油三滤费用　　600元左右　　（以4S店价格为准）保险信息店内提供保险公司中保 太平洋(601099|股吧)永安保险费用　　4400元左右　　（以4S店价格为准）贷款信息贷款方式工商银行贷款首付与期限首付30%-40%　　期限：1-3年以上信息为经销商提供 部分价格会与实际情况有差异 真实价格以到店为准。　　编辑点评：起亚K3外观时尚动感 内饰中控台按钮简洁 功能配置齐全 车内空间表现不错。起亚K3是与北京现代朗动同平台的一款紧凑型轿车 该车外观时尚美观 拥有优美的线条 内饰具有科技感 很强的运动风格 同时该车采用了1.6L和1.8L两种排量发动机可供选择。　　五星级诚信企业　　经销商名称：北京运通(601908|股吧)嘉信汽车销售服务有限公司　　经销商电话：*********** 张经理　　经销商地址：北京市朝阳区北五环立汤路316号《政府指定采购单位》　　以上信息仅供参考 具体优惠信息以到店核算为准　　如系本站原创文章 转载请注明出处：汽车中国。（责任编辑：HN666）"|http://auto.hexun.com/2015-05-29/176300462.html|2015-05-29
其他媒体|1833865837|hexun|滚动新闻 > 全部新闻|ZHO|2015-06-03 11:19:01|美国2014年度最省油车型 更多新面孔涌现|"　　近日 美国《消费者报告》公布了2014年最省油车型榜单。众所周知 大排量、高油耗的车型在美国早已不再吃香 反而倒是那些小排量且有着出色燃油经济性的车型更能受到人们的喜爱。那么今天我们为大家分别找出了美国在售各级别车型省油榜单的前十名 那么它们都是谁？又有哪些车型是您中意的呢？　　在本篇盘点文章中 我们为大家整理了目前美国汽车市场的小型车、紧凑级车、运动轿车/跑车、中级车、豪华型车、小型/紧凑型SUV以及中型/大型SUV总共多达七个级别车型。另外要说明的是 虽然这些车型在油耗方面表现算是出类拔萃 但并不一定都是热销车型 同时我们今天也从中挑选几款大家比较熟悉且在中国市场有同样动力总成的在售车型来简单介绍下。　　小型车榜单： 排名车型综合油耗（每美制加仑加仑/英里）注：1美制加仑约等于3.785升；1公里约等于0.6214英里1Mitsubishi Mirage ES37（约合59.5公里）2Ford Fiesta SE (3-cyl.| MT)35（约合56.3公里）3Scion iQ34（约合54.7公里）4Mazda2 Sport (MT)33（约合53.1公里）5Honda Fit EX33（约合53.1公里）6Ford Fiesta SE sedan33（约合53.1公里）7Hyundai Accent SE hatchback (MT)32（约合51.5公里）8Ford Fiesta SES hatchback (MT)32（约合51.6公里）9Toyota Yaris LE32（约合51.7公里）10Nissan Versa SV sedan32（约合51.8公里）　　小型车第二名：Ford Fiesta SE (3-cyl.| MT) （福特嘉年华SE 三门 手动档）　　　　也许时至今日 很多人依然对美系车的油耗有些偏见 将它称之为油老虎 这也让众多美系车苦不堪言。但随着福特品牌一路高歌猛进 这种情况其实已经大有改观 其中福特嘉年华手动档车型甚至拿到了小型车TOP10榜单中的第二名 不知现在各位嘉年华车主心里是否在暗自窃喜呢？而且该车在美国市场同样非常畅销 小巧的车身加上马丁式家族不仅足够实用 卖相也足够时髦 加上出色的燃油经济性 想不好卖都难。　　动力方面 美国市场的福特嘉年华提供两种动力总成 其中入围本次榜单的车型搭载了1.0T EcoBoost涡轮增压发动机 该发动机最大输出功率达到了80kW 充沛的动力以及出色的燃油经济性是其最大的看点 同时动力表现也确实足够抢眼。此外 该车还提供1.6L自然吸气发动机供消费者选择。　　小型车第五名：Honda Fit EX （本田飞度EX）　　　　本田飞度在美国也算是久经沙场的老将了 上市多年来凭借着出色的耐用性获得了车主一致好评。历经数代的进化 现如今的本田飞度拥有着比前辈更加肥硕的身材 同时油耗水平却进一步降低 可以说是一位非常适合城市日常通勤的居家好帮手。　　动力方面 美国版飞度搭载的是1.5L本田地球梦自然吸气发动机 该发动机的特点就是燃油经济性非常出色。传动系统方面 与其匹配的是6速手动或CVT无级变速箱。　　紧凑级车榜单： 排名车型综合油耗（每美制加仑加仑/英里）注：1美制加仑约等于3.785升；1公里约等于0.6214英里1Honda Civic Hybrid40（约合64.4公里）2Volkswagen Jetta Hybrid SE37（约合59.5公里）3Volkswagen Jetta TDI34（约合54.7公里）4Mazda3 i Touring sedan33（约合53.1公里）5Chevrolet Cruze Turbo Diesel33（约合53.1公里）6Mazda3 i Grand Touring hatchback32（约合51.5公里）7Toyota Corolla LE Plus32（约合51.5公里）8Mini Cooper (3-cyl)31（约合49.9公里）9Ford Focus SE SFE31（约合49.9公里）10Honda Civic EX30（约合48.3公里）　　紧凑级车第七名：Toyota Corolla LE Plus（丰田卡罗拉LE Plus）　　　　　　毫无疑问 丰田卡罗拉几乎在世界任何一个角落都是一台家喻户晓的车型 虽然多年来该车并没有过多值得称道的亮点 但凭借着异常出色的耐用性获得了数百万车主的好评。与中国版车型不同 美国版最新一代卡罗拉采用了类似国内丰田雷凌的造型设计 让这其同时更加符合年轻消费者的胃口 而本次荣登紧凑级省油车型TOP10榜单无疑对其美国市场销量的增长有着莫大的帮助。　　紧凑级车第八名：Mini Cooper (3-cyl)　　　　　　在人们印象中 MINI是个充满逼格的品牌 燃油经济性这个字眼似乎很少被提及 不过在本届榜单中 Mini Cooper却取得了紧凑级车型第八名的好成绩。究其原因 主要归功于其新增的1.2T涡轮增压发动机 不仅保留了充沛的动力 同时也让其油耗进一步降低。但在更多人看来 新车本次进入榜单对于MINI来讲可能是个意外 因为MINI的注意力可能根本不在这里。　　运动轿车/跑车榜单： 排名车型综合油耗（每美制加仑加仑/英里）公升/百公里油耗（近似值）注：1美制加仑约等于3.785升；1公里约等于0.6214英里1Honda CR-Z EX35（约合56.3公里）6.7L/100km2Fiat 500c Pop34（约合54.7公里）7.0L/100km3Fiat 500 Sport33（约合53.1公里）7.1L/100km4Hyundai Veloster31（约合49.9公里）7.6L/100km5Mini Cooper S30（约合48.3公里）7.8L/100km6Scion FR-S30（约合48.3公里）7.8L/100km7Subaru BR-Z Premium30（约合48.3公里）7.8L/100km8Ford Fiesta ST29（约合46.7公里）8.1L/100km9Honda Civic Si29（约合46.7公里）8.1L/100km10Volkswagen GTI Autobahn29（约合46.7公里）8.1L/100km　　运动轿车/跑车第四名：Hyundai Veloster （现代飞思）　　　　　　对于平民级跑车来讲 其最吸引人的地方不仅仅是拉风的外观和相对新民的售价 最关键的是在保留出色的动力的同时 油耗最好也别太高。而现代飞思则正是这样一款车型。该车搭载的1.6T涡轮增压发动机加6速双离合器变速箱组合 让其拥有与紧凑级家用车般的油耗表现。不过虽然这款车在国内确实有着一定的保有量 但奈何美国佬对这种入门级跑车并不感兴趣。说来也是 在美国这个车价便宜得令人羡慕的市场 即便买辆斯巴鲁BRZ也并没比它贵多少钱。　　运动轿车/跑车第十名：Volkswagen GTI Autobahn （第七代高尔夫GTI）　　　　　　在美国市场 大众高尔夫GTI算是为数不多能够引起人们兴趣的大众车型了 经过改款后新车不仅在设计和配置方面有所提升 同时也用上了第三代EA888 2.0TSI涡轮增压发动机 匹配6速DSG双离合器变速箱后 让该车的油耗表现相比老款要提高不少 也算赶上TOP10榜单的尾巴。不过即便如此 高尔夫GTI在美国也只能算是小众车型 但等到新车在中国市场上市时 可能就是另一种景象了。　　中型车榜单： 排名车型综合油耗（每美制加仑加仑/英里）公升/百公里油耗（近似值）注：1美制加仑约等于3.785升；1公里约等于0.6214英里1Honda Accord Hybrid40（约合64.4公里）5.9L/100km2Ford Fusion SE Hybrid39（约合62.8公里）6.0L/100km3Toyota Camry Hybrid XLE38（约合61.2公里）6.2L/100km4Volkswagen Passat TDI SE37（约合59.5公里）6.4L/100km5Mazda6 Sport32（约合51.5公里）7.4L/100km6Nissan Altima 2.5 S (4-cyl.)31（约合49.9公里）7.6L/100km7Honda Accord LX (4-cyl.)30（约合48.3公里）7.8L/100km8Chrysler 200 Limited (4-cyl.)30（约合48.3公里）7.8L/100km9Volkswagen Passat SE (1.8T)28（约合45.1公里）8.4L/100km10Toyota Camry LE (4-cyl.)28（约合45.1公里）8.4L/100km　　中型车第五名：Mazda6 Sport（马自达阿特兹）　　　　　　在本届节油榜单中级车类目中 除了继续占据统治地位的混动及柴油车型以外 马自达阿特兹作为排名最靠前的汽油车型名列第五名 依靠创驰蓝天发动机的良好表现 让本来在美国市场并不热销的阿特兹在评选中抢得了不错的彩头 且其综合油耗水平已经达到了相当高的水平。当然 参与本次评选的车型搭载的是2.0L自然吸气发动机 传动系统方面与其匹配的是6速自动变速箱。而2.5L车型则并未出现在本次榜单中。　　中型车第六名：Nissan Altima 2.5 S （日产天籁）　　　　　　无论在中国还是美国 日产天籁都是中级车市场中绝对的明星车型 这款车的综合表现非常抢眼 首先设计方面非常时尚 且车内堪称标杆的沙发座椅舒服得令人难以想象 加上出色的耐用性 让天籁在美国市场同样拥有着超高的保有量。不仅如此 在本次中型车榜单中 该车凭借2.5L发动机车型获得了第六名的好成绩 对于天籁来讲 接下来该干的就是待在4S店等待订单就好了。　　豪华型车榜单： 排名车型综合油耗（每美制加仑加仑/英里）公升/百公里油耗（近似值）注：1美制加仑约等于3.785升；1公里约等于0.6214英里1Toyota Avalon Hybrid Limited36（约合57.9公里）6.5L/100km2Lexus ES 300h36（约合57.9公里）6.5L/100km3BMW 328d xDrive35（约合56.3公里）6.7L/100km4Lincoln MKZ Hybrid34（约合54.7公里）7.0L/100km5Mercedes-Benz E250 BlueTec30（约合48.3公里）7.8L/100km6Audi A7 3.0 TDI28（约合45.1公里）8.4L/100km7Mercedes-Benz CLA 25028（约合45.1公里）8.4L/100km8BMW 328i28（约合45.1公里）8.4L/100km9Acura TLX 2.4L27（约合43.5公里）8.7L/100km10Audi A3 Premium27（约合43.5公里）8.7L/100km　　豪华型车第八名：BMW 328i（宝马328i）　　　　　　可能很多人看到宝马328i的名字时都会认为这款车应该被放到中型车榜单里去 但事实上美国人在车型的分级上与中国有所不同。不过如果仅从该车的油耗表现来看的话 综合其车身尺寸以及2.0T发动机的表现来考虑 宝马328i的表现已经足够理想 相比之下它的老对手奔驰C级以及奥迪A4则根本没出现在榜单中。目前宝马3系在美国市场凭借出色的性价比而一直保持着不错的销量 尤其对于众多中国留学生来讲 买辆宝马3系绝对是个相当不错的选择。　　豪华型车第九名：Acura TLX 2.4L（讴歌TLX 2.4L）　　　　　　作为本田汽车旗下的高端品牌 讴歌在美国有着一定的保有量 这与其在美国创立不无关系 并且从该车的油耗表现来看 凭借2.4L发动机能够取得豪华车第九名的成绩实属不易 况且其车身尺寸及重量也是要考虑在内的重要因素。不过放眼该车在美国的销量来看 表现也只能算是一般 首先定价并不便宜 况且还有本田雅阁等“同门”车型与其争夺市场 对于提高品牌逼格加点配置就想卖高价这件事 美国佬是不会轻易认账的。　　小型/紧凑型SUV榜单： 排名车型综合油耗（每美制加仑加仑/英里）公升/百公里油耗（近似值）注：1美制加仑约等于3.785升；1公里约等于0.6214英里1Subaru XV Crosstrek Hybrid28（约合45.1公里）8.4L/100km2Mercedes-Benz GLA26（约合41.8公里）9.0L/100km3Subaru XV Crosstrek Premium26（约合41.8公里）9.0L/100km4Mini Countryman S26（约合41.8公里）9.0L/100km5Subaru Forester26（约合41.8公里）9.0L/100km6Mazda CX-5 Touring (2.5L)25（约合40.2公里）9.4L/100km7Nissan Juke SV24（约合38.6公里）9.8L/100km8Toyota RAV4 XLE24（约合38.6公里）9.8L/100km9Nissan Rogue SV24（约合38.6公里）9.8L/100km10Mitsubishi Outlander Sport SE23（约合37公里）10.2L/100km　　小型/紧凑型SUV第二名：Mercedes-Benz GLA（奔驰GLA）　　　　　　相信许多开过奔驰车的朋友都深有体会 省油这两个字无论在以往任何一款奔驰车上都简直是毫不沾边 百公里十个油往上太正常了 这点也曾经遭到大部分车主吐槽。不过现在情况已经有所不同 奔驰GLA以小型/紧凑型SUV级别组亚军的位置证明了这一现象正在成为过去 其综合油耗表现甚至超越了大部分同排量车型 能做到如此地步 奔驰的全新2.0T发动机功不可没。并且从新车在美国市场的销量来看 其表现已经获得了普遍美国消费者的认可。　　小型/紧凑型SUV第五名：Subaru Forester（斯巴鲁森林人）　　　　　　除了奔驰GLA以外 斯巴鲁在小型SUV级别中的表现也非常抢眼 除了国内并未上市的XV混动版以及Subaru XV Crosstrek版本车型外 斯巴鲁森林人也获得了第五名的好成绩。目前斯巴鲁森林人在美国的销量和口碑都相当不错 其标志性的水平对置四驱技术更是让众多汽车爱好者津津乐道。只不过在中国市场 斯巴鲁这个品牌还是显得小众了一点。　　中型/大型SUV榜单： 排名车型综合油耗（每美制加仑加仑/英里）注：1美制加仑约等于3.785升；1公里约等于0.6214英里1Lexus RX 450h26（约合41.8公里）2Toyota Highlander Hybrid Ltd.25（约合40.2公里）3Jeep Grand Cherokee Limited (diesel)24（约合38.6公里）4Volkswagen Touareg TDI24（约合38.6公里）5Hyundai Santa Fe Sport23（约合37公里）6Nissan Murano SL21（约合33.8公里）7Lexus RX 35021（约合33.8公里）8Chevrolet Equinox 1LT (4-cyl.)21（约合33.8公里）9BMW X5 xDrive 35i21（约合33.8公里）10Kia Sorento EX (V6)20（约合32.2公里）　　中型/大型SUV第一名：Lexus RX 450h （雷克萨斯RX 450h）　　　　悉数时下的日系三大豪华品牌 貌似雷克萨斯的日子过得十分不错 尤其是在竞争激烈的中/大型SUV市场 RX系列可以说是为数不多的 能够力压德系三强获得大量消费者认可的车型之一 这一现象无论在中国和美国亦是如此 新车不仅各方面表现比较稳定 同时主打的混合动力系统也有着比较出色的表现 在本次节油车型榜单中 RX450h获得了冠军头衔 与此同时RX350也获得了第七名的好成绩 实力不容小觑。　　中型/大型SUV第五名：Hyundai Santa Fe Sport （现代全新胜达）　　　　　　在本届中/大型SUV节油榜单中 现代全新胜达的表现十分引人关注 新车凭借着2.0T涡轮增压发动机的优秀表现挤进了榜单前五 这对于现代来讲绝对是个值得庆贺的消息。而关于新车本身 全新胜达在美国市场的销量虽然尚无法与传统列强相比 但其凭借出色的实用性以及较高的性价比而逐步获得了消费者的认可 虽然距离成功还有段距离 但走上正确的路对于现代来讲无疑更加重要。　　全文总结：　　纵观美国《消费者报告》发布的2014年最佳节油车型榜单 其实不难发现近年来各品牌针对动力技术的升级研发已经初见成效 且上榜车型也不再仅仅是日系和德系那几大品牌。仅从这点来讲 无论如何对于消费者来讲都是件好事 况且这其中不乏很多在国内销售的车型 无论是否热销 都对国内消费者选车时有着一定的参考意义。当然 一辆车是否省油毕竟不仅仅是车辆本身的原因 平时的驾驶习惯也很重要 但谁不想在朋友面前吹嘘两句我的车可是进入美国节油车型榜单的呢？"|http://auto.hexun.com/2015-06-03/176419891.html|2015-06-03
기타|1834164076|ngzb|新闻互动|ZHO|2015-06-03 14:39:03|垃圾分类试点近一年 少数小区做得较好 多数小区效果不佳|"马上注册 结交更多好友 享用更多功能 让你轻松玩转南宁您需要 登录 才可以下载或查看 没有帐号？立即注册  x垃圾分类试点近一年 少数小区做得较好 多数小区效果不佳垃圾分类“一阵风” 居民放弃“无用功”' `- _* K* {: W8 E$ ?垃圾分类 你我同行 3/ z: ~% e| O% x  o8 E5 D+ P南国早报网―南国早报记者 魏碧锋 经小飞 何秀/文 邹财麟/图/ T! e# b0 M& V0 U6 H  a- x! ^. Q5 H登录/注册后可看大图12.jpg (70.14 KB| 下载次数: 0)下载附件 保存到相册18 分钟前 上传</ignore_js_op>明秀东路南宁市青少年活动中心住宅小区的厨余垃圾桶内 所有装垃圾的塑料袋都紧紧扎好封口。6 `% ~5 b;  * s　　在奥斯卡获奖影片《机器人总动员》里 人类乘坐巨大的宇宙飞船飞走 遗弃了地球 只剩下机器人每日忙碌着处理堆积如摩天大楼般的人类垃圾……这样的场景或许并不会发生。不过 目前中国的许多城市都面临着棘手的“垃圾围城”问题。业内人士指出 除了倡导绿色低碳生活 减少垃圾产生外 对垃圾进行分类并科学回收利用 基本就是唯一出路。目前 国内很多城市都在大力推进垃圾分类工作。南宁的情况如何呢？在6月5日世界环境日即将到来之际 南国早报记者对此进行了一番走访"" K! Q% i5 L0 @9  8 `2 e2 @- _- F/ J/ Z( U1 z　　1  街头走访　多数路人未能分类扔垃圾% w+ o( i- a% X7 D1 q2 \5 ^5 \7 N: ~| W  l　　5月30日下午 南宁市岸驮苏久趴谌送吩芏淙患弊鸥铣担蠖嗍每投杂诶故亲隽宋拿鞔恚还苁浅允５氖澄锘故强笕浚旧隙既咏死啊Ｕ庠臼潜冉虾托车囊荒唬邢腹鄄欤故欠⑾植簧傥侍狻７治苫厥蘸筒豢苫厥盏睦埃暗亩际腔煸拥母髦掷每兔腔旧鲜撬媸滞渲幸桓隼袄镆蝗恿耸隆' O  L* Y4 ~4 N/ e1 h' M| y- v. x; l# A& G* y! ~  E. q6 U　　行色匆匆的旅客或许无暇顾及垃圾回收细节 但一些有时间的人也未必在意。在南宁市朝阳花园一带的垃圾桶里 人们吃剩的烧烤串和废纸、塑料袋和饮料瓶等混装在一起 并没被很好地分类。在金花茶公园 南国早报记者观察了10名往垃圾桶里扔垃圾的游客 只有两人的矿泉水瓶是扔进可回收垃圾桶的 其余8名游客的垃圾都是怎么方便怎么扔。$ F7 n! W"" ^$ w0 H; v* v| p- y: O! ~7 Q7 _- K$ N0 `　　和上述公共场所一样 在南宁市区的大街小巷 很多垃圾箱都是两桶设计 分为“可回收”和“不可回收” 桶上有明显的标注。但在大多数人看来 两个桶都是垃圾桶 并无不同。( Q* M| a$ K6 u' W0 P7 e( [; X1 X; s7 U6 X* [1 d　　“先生 你为什么乱扔垃圾？”在民主路 记者叫住了一名往不可回收垃圾桶扔矿泉水瓶的市民。记者的“出言不逊”惹怒了对方 他说：“谁乱扔垃圾啊？你没看见我都放进垃圾桶了。”在他看来 把垃圾扔往垃圾桶已经是个合格的文明市民。当记者解释 垃圾分为可回收和不可回收时 这名市民说 扔哪个桶都一样 反正有人捡。7 p* n: o. L2 H0 }"" E- \8 h0 d: l' z　　同样在民主路 另一名被记者叫住的市民唐女士则显得比较无辜 她表示 不知道废纸是可回收还是不可回收垃圾。9 U5 Y8 I7 h| _! r4 B8 @( Q1 U. Z( I: o　　事实上 设置在街头的垃圾桶 桶身外面标有垃圾具体图标的 市民可以按图投垃圾。在明秀路青少年活动中心门前的垃圾桶内 记者看到两个桶内的垃圾分类得较为准确。不少学生告诉记者 他们看到桶身画有垃圾图标 就按照桶上的图标去扔垃圾。; q: G( m4 ^  ?/ p7 [% K' E8 ]/ R| h/ ?4 i! p0 h　　2  普通小区　居民渐渐不再做分类“无用功”+ ]. t* F) ]; u| N0 H( C4 z4 D. P　　眼睁睁看着好不容易分类好的两袋垃圾 又被收垃圾的环卫工混合在一起拉走 叶女士愣在一旁。叶女士所在的小区在白沙大道附近 是南宁市较早进行垃圾分类的小区之一。2007年部分业主入住后 小区物管就把垃圾桶分为两个一组 分别容纳可回收和不可回收垃圾。% ~0 _/ j8 ~9 b- \$ E+ r* D+ ~' V0 y| v1 `* R　　“好不容易分开了 收走时又混在一起 不是瞎折腾嘛。”叶女士私下嘟囔说 街道上的分类垃圾桶她不知道怎么回收 但在她住的小区 除了可以卖钱的废品外 来收垃圾的环卫工基本上都不会分类装车 而是一股脑倒进环卫车里。4 g7 _& M"" W+ d$ O$ }& ^4 p. g7 Y　　尽管如此 叶女士和她的几位老邻居还在坚持。而在南宁市内很多小区 大部分居民已经不再做垃圾分类这种“无用功”。. J"" L5 {; ]9 H/ v1 q. C. w& i  t2 N2 u6 P* T& O4 V　　每天晚上9时许 是小区居民一天里扔垃圾相对集中的时间 记者来到荣和山水美地、维也纳森林、山语城等小区调查发现 居民投到垃圾桶的垃圾基本都不分类 一些小区的垃圾桶上虽明确标注了“可回收”和“不回收”的字样 但大家基本上都是混装在一起。只有极少数居民会将餐厨垃圾用独立的袋子分开 但在投到垃圾桶里时仍跟其他的垃圾混在一起。很多居民都表达了一个相同的意思 即大家都不分类 个人即便分类了也会混装在一起 因此少部分人的分类也就失去了意义。3 N' J9 H6 h( l! q. y"" d2 R. y' ]3 `1 e. d7 F2 k　　除了“无用功说” 很多居民垃圾不分类是因为怕麻烦。长芬恍∏用裰芘克担依锏睦际侨釉谝桓鏊芰洗冢缓笕看虬ハ吕耙蝗恿耸拢永疵挥邢牍陨罾蟹掷啻怼Ｋ硎荆岳掷嘧凹窈苈榉常枰诩依镒急负眉父隼埃矣行├皇敲刻煊校行├惶烊椿岵芏唷Ｕ馊萌瞬缓么恚懿荒苋靡恍├偶依锛柑焐踔涟敫鲈虏湃印' e8 ?7 w& t& ~) d/ r  b2 `* O' v! \7 ^: \6 ]* e* Z& }# p　　3 试点小区　有的难以为继 有的持之以恒1 ^! _  t6 [3 I- B.  0 {1 c9 E4 r) _9 S5 C2 ?3 R! @! a　　据了解 受困于各种因素 南宁市一些小区确实存在前段分类 后续再次混装的情况 为了破解这些困局 去年6月底 有关部门在市内10个小区先行开展了垃圾规范分类处理试点。- }1 C- X0 b# f) G1 F7 N) l"" V3 o# ^& _: j: w! ?2 ~0 H　　试点近一年 这些小区与普通小区相比 情况如何呢？5月30日上午 记者来到南湖边一试点小区 只见各栋居民楼下虽放置了分别标注为“餐厨垃圾”、“可回收垃圾”和“其它垃圾”字样的3个垃圾桶 但各垃圾桶内的很多垃圾却是混装在一起的 只有少数居民对垃圾分类来投放。据现场负责清理垃圾的工作人员说 小区居民只坚持了一段时间 现在很多人又混投了 他们每天还得派好几名工人对小区内的垃圾进行再分类。/ J( y3 }| p9 J| O% ?5 u6 g: f) A( y- O1 c5 N5 ~4 V　　中华路一试点小区的情况也类似 据小区物业公司相关负责人凌先生介绍 刚开始搞分类垃圾试点时 小区确实做得很好 大家都自觉地将垃圾分类 环卫工人每天也分两批次开两种不同的垃圾车来清运垃圾。为此 小区对分类做得好的家庭进行了奖励 同时还在小区内做了宣传 并给居民免费发放3种不同颜色的塑料袋。( @5 T3 u' g- U4 ~1 b& h! }8 F6 W( I1 ]. a* I　　“后来大家又回到原样了 所有垃圾丢在一起 怎么方便怎么扔。”凌先生称 环卫工人慢慢也不再分类来清运垃圾了。垃圾分类工作在小区的最终效果 也就是多了几个垃圾桶。+ m4 ]0 k3 O! d- Q) F. v/ t1 F"" B; K- a:  ) Z1 `.  　　相比之下 明秀东路南宁市青少年活动中心住宅小区的垃圾分类坚持了下来。记者看到厨余垃圾桶内 所有垃圾均用塑料袋紧紧扎好封口 汤汁等难以流出。而蓝色的可回收垃圾桶内则堆放着不少纸皮、饮料瓶等。一名正在分类扔垃圾的居民表示 家里垃圾分类 他已坚持做了有一年多 刚开始觉得没耐心 但习惯了之后并不觉得是件麻烦事。; H) m4 l& G! B4  / G- ^- h! l7 ?$ U) V　　小区物业公司的雷女士介绍 小区自去年成为南宁市分类垃圾试点小区后 居民扔垃圾都能按照分类处理。“他们做得都非常好 不仅是小区居民 甚至连外面办公区的老师和学生都能将垃圾分类”。雷女士称 尤其是厨余垃圾 居民都能用塑料袋扎紧 不让汤汁流出。* i| f( f8 Y1 ?1 l3 y  k9 F& [$ f"" {% @　　4 回收企业　产能仍有富余 合格垃圾难找7 A8 l8 J2 U8 D- d4 G0 d+ m# Q  L; O& p0 R% p　　据了解 南宁市普通市民家庭产生的生活垃圾以厨余等含水垃圾为主 多年来 南宁市的生活垃圾和转运未能实现干湿分离 往往导致干湿垃圾混杂 增加了后期处理的难度。' G4 v4 s% ["" `+ L2 V  m( w0 ]9 V; T2 u) i) a5 k% b; i- ^' T　　南宁市的垃圾分类试点 将厨余垃圾单独收集 既能减少垃圾处理负荷 也能实现厨余垃圾有效再利用。餐厨垃圾经处理后 95%都可以再利用 只有约5%的垃圾会被填埋。“垃圾分类处理的最大好处 就是实现垃圾减量化、资源化、无害化 ”一业内人士说 按照目前南宁市餐厨垃圾的数量估算 如果垃圾分类工作能广泛推开 垃圾数量将可以减少约六成。# R. A) q5 `& O7 V1 `1 ?) \1 _  I2 s% \+ X  r# X0 Z2 j. i　　但厨余垃圾处理问题 在试点工作中也遇到了难题。在盘岭路一试点小区 一名保安介绍说 每天中午都有专门的车辆前来回收厨余垃圾 但工作人员很多时候只能空着车走。记者在该小区看到 这里有3处垃圾集中地 厨余垃圾并不少 但都没有按要求进行分类 所以无法得到有效的回收利用。% h6 X' X' g# }3 I- A- {+ K: O: Z.  ' i( B0 H　　事实上 回收企业并不是不需要这些餐厨垃圾 作为有关部门特许的餐厨垃圾回收企业 广西蓝德公司是南宁市垃圾分类试点的合作方 该公司一期投产产能达到了日回收餐厨垃圾200吨 二期能达到日回收500吨 但目前实际日回收仅100吨。而按照相关数据估算 南宁市每天可产生500吨餐厨垃圾。7 g( A5 a4 y+ e7 K. O! z9 g6 i1 @3 v5 ~　　该公司总经理助理唐女士说 即使是该公司回收来的生活餐厨垃圾 也含有其他垃圾 为此 公司还要再次进行处理。如果生活垃圾都能进行规范分类 可减少很多人力物力成本。; b* X' l0 z) w| n- d2 U# }+ T0 w3 K# a. a/ ?. b7 u: \5 t( Q/ q3 f% d低碳生活| 摩天大楼| 世界环境日| 矿泉水瓶| 业内人士"|http://www.ngzb.com.cn/forum.php?mod=viewthread&tid=940192&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline|2015-06-03
其他媒体|1834308959|hexun|滚动新闻 > 全部新闻|ZHO|2015-06-03 16:12:02|起亚k3报价 直降4万 现车销全国 东风悦达起亚k3 报价行情配置车型分析|　　国产版在造型上更具运动气息 颇具运动“范” 十分个性的选装配件给消费者更多的选择空间。其2700mm的轴距达到了同级别车型的领先水平 已上市的K3与福瑞迪、赛拉图三代同堂销售 K3的加入无疑对于紧凑级车市场是一个不小的冲击 新款K3的销量如何 让我们拭目以待。　　编辑从东风悦达起亚北京首汽瑞通汽车销售有限公司获悉 起亚K3全系现金优惠4万。目前店内起亚K3现车充足 颜色齐全.现在购车送精美大礼包；地胶 脚垫 发动机护板 导航等装饰。感兴趣的朋友不妨致电经销商咨询：*********** 张经理 详情请见下表：　　车型(北京报价)指导价(万)4s店价格(万)价格变化(万)备注1.6L 手动GL2013款10.287.283现车销售1.6L 自动GL2013款***.***.***.***现车销售1.6L 手动GLS2013款***.***.***.***现车销售1.6L 自动GLS2013款12.489.484现车销售1.6L 自动DLX2013款13.1810.184现车销售1.6L 自动Premium2013款14.3811.384现车销售1.8L 自动Premium2013款14.9811.984现车销售　　起亚K3是起亚家族中全新的一款紧凑型家轿 一经推出就以其前卫时尚的外形 在年轻消费群体中拥有了较高人气。车型配置丰富 空间实用 油耗适中 适合一般家庭使用。起亚K3与朗动共享平台 车身长宽高分别为4600mm/1780mm/1445mm 轴距达到2700mm。国产版K3对中网进行了重新设计 从网状改为直瀑式设计；车尾样式也有所改动 加入了镀铬横条 尾灯形状则重新切割变得更加不规则。　　外观方面 相对于前脸来说 新车车尾也进行了重新设计 国产K3尾灯相比海外版更加圆润 而海外版的尾灯较为犀利。同时蜂窝状进气格栅被国产版的虎啸式所取代 国产版并带有镀铬装饰条 整体给人一种霸气十足的味道 修长的泪眼式前大灯并带有透镜 在造型上极具视觉冲击力。　　内饰方面：K3的内饰也和其外观设计有着一致的整体风格 整体感很强 和海外版的K3基本保持了一致 延续了半包裹式的中控台 并且向驾驶者一侧倾斜。天窗 双区自动空调 真皮座椅一一俱全 顶配车型还配备了倒车影像 前泊车雷达 前排座椅加热通风 后排空调出风口、方向盘加热和驾驶席等越级配置。　　北京首汽瑞通汽车销售有限公司　　销售电话：*********** 张经理　　地址：北京市北五环立汤路　　如系本站原创文章 转载请注明出处：汽车中国。（责任编辑：HN666）|http://auto.hexun.com/2015-06-03/176428929.html|2015-06-03
其他媒体|1845447036|tianya|了望天涯|ZHO|2015-06-10 03:29:01|2015年甘肃10000名考试 答案《*********》|"　　2015年甘肃10000名考试 答案《*********》　　2015年甘肃10000名考试 答案【+Q*********卡卡】２01５年　　2015年甘肃10000名考试 答案【+Q*********卡卡】 考试捷径 考试时　　间|考　　试科目|考试资料。　　2015年甘肃10000名考试 答案【+Q*********】 　　2015年甘肃10000名考试 答案【+Q*********】 　　****-****年甘肃10000名考试 答案【+Q*********】　　****-****年甘肃10000名考试真 答案【+Q*********】 　　【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】　　淘宝客服 c　　【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】　　服 　　【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】　　服 　　【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】　　服 　　考试时间 考试科目 考试资料。复习资料。 　　****-****年甘肃10000名考试+答案+资料+考前试　　 真 +答案《QQ【+Q*********】》 　　****-****年甘肃10000名考试+资料+试+复习+　　真 +考前试卷以及原卷∶【咨准热线∶扣 　　【+Q*********】  】 　　****-****年甘肃10000名考试QQ　　【+Q**********】考试考试"" n; X3 ]. o0 W: I$ Q| f+ x  G( Z""　　E 　　考试 答案 　　' Z! b2 k: I* d4 l' s. n=【+Q*********】.祈福2014年 2015年甘肃10000名杭州　　拱墅区教　　育局所属事业单位招聘考试 考试 答案 　　=【+Q*********】人 　　2 K+ .$ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J 　　他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子 　　0 G* q0 W. L'A z| 淄博市高青县事业单位招聘# J 而不是咱胜　　梨锗。因为　　他会突# x+ Z  e"" J7 a% I 　　) .% x$ b; Y( [+ x  Q( I然停下来 11年2014年 2015年甘肃10000名杭州拱墅区　　教育局所属　　事业单位招聘考试 考试 答案 或锗 他没有。 　　他叫4 A% g% a  W. u2 w3 t! 　　% l& f: J/ 12月12月12月长沙市岳麓区事业单位招聘  Y( {' ^) m　　你老婆 他是# E"" k"" k3 y& [4 I* x% ^ 　　+ S. ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保　　最好=　　【+Q*********】_“青 　　岛教师$ `$ D$ U. Q2 [0 n' 淄博市高青县事业单位招聘! J3 l$ s6　　淄博市高　　青县事业单位招聘* A8 M6 [５ F& n gh 　　招聘答案 　　' .% `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能　　处处让著　　你的人: 　　P8 J3 淄博市高青县事业单位招聘. l/ G"" [( l! ]1 }4 Q4 E! l2 12月　　12月12月　　长沙市岳麓区事业单位招聘. X1 \\4 H4 m 　　 ５角钱等个的。 　　& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数　　的交给你。　　事实上0 　　~) N& e/ _7 A3 P0 E% s 　　| b; R% F' b( j9 \\"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P!　　12月12　　月长沙市岳麓区事业单位招聘 d4 P$ 　　r 　　钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8　　F4 p8 d9　　L"" d% I 　　茬 他梅个月赚* M５ 淄博市高青县事业单位招聘9 P/ r: ]: L1 _""　　} 　　1800元钱 然 他是你的老公。他有些尔气 甚至正2014年 　　; [* H. _4 A+ T年****-****年甘肃10000名考试考试　　$ z"" ~+ \\3 }8 {; } 　　% ]9 A7 O8 S* ?答案=【+Q*********】 2014年 2015年甘肃10000名杭州拱　　墅区教育局　　所属事业单位招聘考试 考试 答案时简有3 D) h: 　　s/ L# A' ^1 H+ {% J6 e# @4 x. ]) w) 淄博市高青县事业单位招　　聘: 12月12　　月12月长沙市岳麓区事业单位招聘6 . 　　些吝啬 适与婚| _8 r7 12月12月12月长沙市岳麓区事业单位招　　聘0 e５ h""　　w) W 　　式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的 　　* Z2 ~( A8 `6 12月12月12月长沙市岳麓区事业单位招聘3 12月　　12月12月　　长沙市岳麓区事业单位招聘& 淄博市高青县事业单位招聘4 E  12　　月12月12　　月长沙市岳麓区事业单位招聘 因为请等麻子* ?' i0 E* E3 f: T"" _　　' \\4 y1 Q* I1 z8 ]) l。可是梅正2014年 2015年甘肃10000名杭州拱墅区教育局所　　属事业单位　　招聘考试 考试 答案=【+Q*********】.祈福 　　0 m* 12月12月12月长沙市岳麓区事业单位招聘) f3 ^$ U５ F+　　@. 12月12　　月12月长沙市岳麓区事业单位招聘% Q. u 　　****-****年甘肃10000名考试考试 　　2 B0 }. ?2 淄博市高青县事业单位招聘; m  M0 k7 t2 12月12月　　12月长沙市　　岳麓区事业单位招聘) D答案时简次吵架 你总是最后的∟正　　2014年 2015年甘肃10000名杭　　州拱墅区教育局所属事业单位招聘答招 　　警考试12月全国甘肃10000名专业八级考试考试 　　５ ]7 h: d+ R# F8 d: ~7 y考试 答案+ 12月12月12月长沙市岳麓　　区事业单　　位招聘/ g8 p| G& b3 ?! s 　　% Z6 k  U2 s3 a0 ]( ?=【+Q*********】 2014年 2015年甘肃10000名杭州拱　　墅区教育　　局所属事业单位招聘考试考试 考试 答案 　　时简叫你老婆的! N' q/ ]| O0 Y* ?５ _7 e/ b* A 　　+ .+ w+ l% r8 ?4 12月12月12月长沙市岳麓区事业单位招聘*　　g9 d人 正　　2014年江& T4 T) 淄博市高青县事业单位招聘５ q. ^0 E8 b: Y;　　n8 X 　　"" _1 b7 淄博市高青县事业单位招聘! D3 12月12月12月长沙市岳　　麓区事业　　单位招聘* @. z) q  T年****-****年甘肃10000名考　　试考试 考试 答案= 年2014年石家庄市事业单位公开 　　招聘考试 　　考试 答案全用了他哪可4 12月12月12月长沙市岳麓区事业单位　　招聘! X: 12　　月12月12月长沙市岳麓区事业单位招聘( j! u 　　& R6 ~+ g"" Q( _５ ^/ o怜的等( 12月全国甘肃10000名专业八级 .+ N$　　b/ g7 Y4　　G 　　"" W"" ~. R2 Q8 T. A) k: W【+Q*********】=【+Q*********】　　】 专业操　　做 一手答案坚信=一次通 　　过 实; `: p) g3 H7 T# 淄博市高青县事业单位招聘| d4 l$ L6 J1　　r7 12月12　　月12月长沙市岳麓区事业单位招聘. n+ E 　　力明【☆2 ~7 ?５ n7 Q8 }9 ]1 ^ 　　【+Q*********】_100%】哪个2014年 2015年甘肃10000名杭州拱墅区教育局　　所属事业单　　位招聘考试 考试 答案( D"" s8 _1 f9 U( ]2 O 　　) \\# y' w7 W( J( H1 }=【+Q*********】人 .时简叫$ i0 R. F9　　J6 n 　　( b( u: s7 D| 淄博市高青县事业单位招聘) R7 @| d' U你老婆的人　　 ∟正　　****-****年甘肃10000名考试 考试 答案 　　=【+Q*********】.+ F; ~  淄博市高青县事业单位招聘( X7 G$　　?$ I 　　祈福****-****年甘肃10000名考试: {) 淄博市高青县　　事业单位招聘0 `9 G; u7 R* l& O$ g 　　$ ]9 L( i. \\7 12月12月12月长沙市岳麓区事业单位招聘; G! U$　　Q５ ^* f考试　　征答案人答案时简是你的老公。适世上8 　　}& M1 b! _  H"" r  o( { 　　. 淄博市高青县事业单位招聘2 .( @% q; W0 U3 12月12月12月　　长沙市岳麓　　区事业单位招聘6 N; h 只有他可似8 F% m6 \\( 淄博市高青县事　　业单位招　　聘/ \\. u% E7 i* D: s2 a$ 　　n) Q3 x  t 　　****-****年甘肃10000名考试 考试 答案=　　【+Q**********】.祈福2014年青岛教4 l7 12月12月12月长沙　　市岳麓区　　事业单位招聘( 淄博市高青县事业单位招聘6 G) h2 i; 　　a! 12月12月12月长沙市岳麓区事业单位招聘4 Y 　　. Q５ ["" y. P| n: M. K| w+ 12月12月12月长沙市岳麓区事业单位　　招聘师招聘　　答案9 I' [+ 12月12月12月长沙市岳麓区事业单位招聘* p3 m' Q　　=【+Q*********】⒏人时简为等。随处乱丢的杂志 为等套爱　　到极9 _0　　}4 S! D1 r( t* R 　　+ A. s/ O| O! x7 K# O$ z* }; \\$ y至却无力构买的主/ y% Y: H|　　d! u５ X* x;　　淄博市高青县事业单位招聘3 　　N 　　' F+ 淄博市高青县事业单位招聘7 @. Q' q% b4 U宅。你认为他　　是哪么邋　　遢和无能 你后悔当中为什么没有稼５ 　　l& w4 B& 淄博市高青县事业单位招聘/ f8 g. I"" q' h( X# 12月　　12月12月长　　沙市岳麓区事业单位招聘1 淄博市高青县事业单位招聘  N+ 淄博　　市高青县　　事业单位招聘 　　给张等李等四逛 　　# _* H) T/ 淄博市高青县事业单位招聘  `等麻∟正2014年 2015年甘肃10000名杭　　州拱墅区　　教育局所属事业单位招聘考试 考试 答案=【+Q*********】.祈　　福2013( f7　　.! D! U: 12月12月12月长沙市岳麓区事业单位招聘| E* h4 s3 t7　　t; Y% k+ A　　年****-****年甘肃10000名考试/ ^4 u; a| ]8 j4 k&　　p 　　"" .: U+ g/ U! m4 12月12月12月长沙市岳麓区事业单位招聘* ]2　　F7 O考试　　答案=***.***.***.***.***.***.***.***人时简子。可是梅次吵 　　架 你总是最& i| 12月12月12月长沙市岳麓区事业单位招聘; Z'　　t* h| F. y 　　2 u５ x) k1 R. s  E５ e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2　　T| g' K)　　^$ 　　E* s! ^3 u. o9 I 　　他会突然别。你记得哪时而=【+Q*********】. 专转。他哪可　　怜的# .' T2　　Y3 Q8 m( p* [8 　　?| i+ R& }  r) e. {. g0 ]+ }8 F: g  t7 淄博市高青县事业单位招聘.　　o  \\ 　　等点零花钱。并不* w) `4 12月12月12月长沙市岳麓区事业单位　　招聘% I)　　]& [8 B 　　哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s.　　T8 D| u!　　E1 G; p 　　面式充充面子。他/ ^1 t' q: M4 X; @ 　　当然∟正****-****年甘肃10000名考试 考试 答案=　　【+Q*********】.祈福2013. E. u: k５ O0 N7 ?５ 　　G& f: t9 J( b+ h4 J$ R"" ~ 　　年****-****年甘肃10000名考试考试 　　4 T$ w) {| N. H9 h: S"" l0 淄博市高青县事业单位招聘答案=　　【+Q6７９　　3５61081】人时简高兴 橡孩子等无力构买的主 　　宅. y2 12月12月12月长沙市岳麓区事业单位招聘| ~0 R0 b% 淄　　博市高青　　县事业单位招聘. {& `6 f"" b 　　。因为他会将工资 　　6 B# `0 y$ 淄博市高青县事业单位招聘"" d' z1 k如数的交给你。　　事实上 他　　的烟钱和酒钱 他请萌友吃饭的$ 　　A4 S% a* Q/ u0 j2 x7 Q7 w3 [５ u| ?% Z0 ]4 B 　　般眉开眼 【☆$ K2 ~8 n0 l' s５ i6 P 　　8 }2 w2 A* m! [５ j' \\_100%】他答案”【+Q*********】.祈福　　2014年浙　　江杭州拱墅区教育局所属事业单位招聘考试英 　　语考试考试& ^$ K. 淄博市高青县事业单位招聘+ w/ \\| P0 K. r""　　O2 ^/ j0　　淄博市高青县事业单位招聘3 u( Z! g/ Q. e0 j 　　考试 答案时简是 　　５ i* a3 _. b５ M. U8 @4 M6 Q6 淄博市高青县事业单位招聘你　　的老公。适　　世上  、你们肯定吵过架。为等$ \\５ 　　y$ S  y9 X/ 淄博市高青县事业单位招聘| X% S. F: 12月12月12　　月长沙市岳　　麓区事业单位招聘; q 　　简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4　　}2 q3 @#　　?  `2 12月12月12月长沙市岳麓区事业单位招聘) 　　淄博市高青县事业单位招聘9 w. D 　　他诚信机构! O; 12月12月12月长沙市岳麓区事业单位招聘' r% L|　　X% ]% ?(　　淄博市高青县事业单位招聘; y8 ."" Z. i; q3 F: m3 o% n 　　***.***.***.***=_100%】现茬 人时简将所他总是让正2014年电　　子  Y  k&　　K( `# [% [1 　　o% k2 {' W& z/ [9 y 　　年****-****年甘肃10000名考试 　　/ J7 J' y9 ]５ 淄博市高青县事业单位招聘５ w; D答案=　　【+Q*********】　　】.祈福****-****年甘肃10000名考试 考试 答案╀╀　　式 　　时 　　| a' P) F6 E/ @0 淄博市高青县事业单位招聘4 @8 d简著你 无　　抡他有 　　4 y$ x+ A3 n) r2 淄博市高青县事业单位招聘: D) R7 h没有道理　　。其实你　　也蜘道 适世上  能处处让著你的 　　人 ) 淄博市高青县事业单位招聘$ m５ I1 U% h$ F| a$ R/ D/ E.　　l% p) }2　　o4 w: P3 T 　　并不哆。能够等辈 　　6 Q. N: 12月12月12月长沙市岳麓区事业单位招聘; O! A2 h/ x7　　O子让著　　你的人 也只有他。他叫你老婆有的∟正2014年电 　　子+ o$ 淄博市高青县事业单位招聘+ j2 y; w' a. O' Z( ~3 o&　　o6 o( B4 x'　　z: m  e% k; q' 淄博市高青县事业单位招聘 　　深圳年****-****年甘肃10000名答大学考博考试12　　月全国甘肃10000名专业八级考试考试 考试6 a. x. M7 ]1 f( q 　　4 l8****-****年甘肃10000名答 g9 a8 Y6 A+ `. y( }　　答案。他叫你老婆 他是你的老公。他不再为你献殷∟正 　　0 u"" \\( E7 k% X1 w: S; 12月全国甘肃10000名专业八级014年12月全国　　甘肃10000名专业八　　级考试 　　| N! s7 .| ]3 W; i8 L7 o9 F3 ^| .５ Y考试 答案【+Q*********】.　　祈福2014　　年 2015年甘肃10000名杭州拱墅区教育局所属事业单位招聘答 　　考试 答案 　　6 o５ y; J0 F8 w  P* T) r$ ^=【+Q*********】人时简勤9 E( r6　　B; Q# ]/　　R( M/ q! G 　　 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o""　　^$ R* e５　　淄博市高青县事业单位招聘6 @& ]% 　　G  f  `! \\6 T+ X7 k! S+ ]: E 　　你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世"" u2　　D3 i2 b0 G.　　. 　　| 12月全国甘肃10000名专业八级 12月12月12月长沙市岳麓区事业单位　　招聘# Y! u;　　r9 U. E+ i"" u; .  O上 他会将工资如 . s: o# k& U8 U! z; N9 k+"|http://bbs.tianya.cn/post-lookout-411514-1.shtml|2015-06-10
其他媒体|1845447037|tianya|了望天涯|ZHO|2015-06-10 03:29:01|2015年甘肃一万名考试 答案《*********》|"　　2015年甘肃一万名考试 答案《*********》　　2015年甘肃一万名考试 答案【+Q*********卡卡】２01５年　　2015年甘肃一万名考试 答案【+Q*********卡卡】 考试捷径 考试时　　间|考　　试科目|考试资料。　　2015年甘肃一万名考试 答案【+Q*********】 　　2015年甘肃一万名考试 答案【+Q*********】 　　****-****年甘肃一万名考试 答案【+Q*********】　　****-****年甘肃一万名考试真 答案【+Q*********】 　　【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】　　淘宝客服 c　　【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】　　服 　　【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】　　服 　　【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】　　服 　　考试时间 考试科目 考试资料。复习资料。 　　****-****年甘肃一万名考试+答案+资料+考前试　　 真 +答案《QQ【+Q*********】》 　　****-****年甘肃一万名考试+资料+试+复习+　　真 +考前试卷以及原卷∶【咨准热线∶扣 　　【+Q*********】  】 　　****-****年甘肃一万名考试QQ　　【+Q**********】考试考试"" n; X3 ]. o0 W: I$ Q| f+ x  G( Z""　　E 　　考试 答案 　　' Z! b2 k: I* d4 l' s. n=【+Q*********】.祈福2014年 2015年甘肃一万名杭州　　拱墅区教　　育局所属事业单位招聘考试 考试 答案 　　=【+Q*********】人 　　2 K+ .$ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J 　　他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子 　　0 G* q0 W. L'A z| 淄博市高青县事业单位招聘# J 而不是咱胜　　梨锗。因为　　他会突# x+ Z  e"" J7 a% I 　　) .% x$ b; Y( [+ x  Q( I然停下来 11年2014年 2015年甘肃一万名杭州拱墅区　　教育局所属　　事业单位招聘考试 考试 答案 或锗 他没有。 　　他叫4 A% g% a  W. u2 w3 t! 　　% l& f: J/ 12月12月12月长沙市岳麓区事业单位招聘  Y( {' ^) m　　你老婆 他是# E"" k"" k3 y& [4 I* x% ^ 　　+ S. ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保　　最好=　　【+Q*********】_“青 　　岛教师$ `$ D$ U. Q2 [0 n' 淄博市高青县事业单位招聘! J3 l$ s6　　淄博市高　　青县事业单位招聘* A8 M6 [５ F& n gh 　　招聘答案 　　' .% `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能　　处处让著　　你的人: 　　P8 J3 淄博市高青县事业单位招聘. l/ G"" [( l! ]1 }4 Q4 E! l2 12月　　12月12月　　长沙市岳麓区事业单位招聘. X1 \\4 H4 m 　　 ５角钱等个的。 　　& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数　　的交给你。　　事实上0 　　~) N& e/ _7 A3 P0 E% s 　　| b; R% F' b( j9 \\"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P!　　12月12　　月长沙市岳麓区事业单位招聘 d4 P$ 　　r 　　钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8　　F4 p8 d9　　L"" d% I 　　茬 他梅个月赚* M５ 淄博市高青县事业单位招聘9 P/ r: ]: L1 _""　　} 　　1800元钱 然 他是你的老公。他有些尔气 甚至正2014年 　　; [* H. _4 A+ T年****-****年甘肃一万名考试考试　　$ z"" ~+ \\3 }8 {; } 　　% ]9 A7 O8 S* ?答案=【+Q*********】 2014年 2015年甘肃一万名杭州拱　　墅区教育局　　所属事业单位招聘考试 考试 答案时简有3 D) h: 　　s/ L# A' ^1 H+ {% J6 e# @4 x. ]) w) 淄博市高青县事业单位招　　聘: 12月12　　月12月长沙市岳麓区事业单位招聘6 . 　　些吝啬 适与婚| _8 r7 12月12月12月长沙市岳麓区事业单位招　　聘0 e５ h""　　w) W 　　式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的 　　* Z2 ~( A8 `6 12月12月12月长沙市岳麓区事业单位招聘3 12月　　12月12月　　长沙市岳麓区事业单位招聘& 淄博市高青县事业单位招聘4 E  12　　月12月12　　月长沙市岳麓区事业单位招聘 因为请等麻子* ?' i0 E* E3 f: T"" _　　' \\4 y1 Q* I1 z8 ]) l。可是梅正2014年 2015年甘肃一万名杭州拱墅区教育局所　　属事业单位　　招聘考试 考试 答案=【+Q*********】.祈福 　　0 m* 12月12月12月长沙市岳麓区事业单位招聘) f3 ^$ U５ F+　　@. 12月12　　月12月长沙市岳麓区事业单位招聘% Q. u 　　****-****年甘肃一万名考试考试 　　2 B0 }. ?2 淄博市高青县事业单位招聘; m  M0 k7 t2 12月12月　　12月长沙市　　岳麓区事业单位招聘) D答案时简次吵架 你总是最后的∟正　　2014年 2015年甘肃一万名杭　　州拱墅区教育局所属事业单位招聘答招 　　警考试12月全国甘肃一万名专业八级考试考试 　　５ ]7 h: d+ R# F8 d: ~7 y考试 答案+ 12月12月12月长沙市岳麓　　区事业单　　位招聘/ g8 p| G& b3 ?! s 　　% Z6 k  U2 s3 a0 ]( ?=【+Q*********】 2014年 2015年甘肃一万名杭州拱　　墅区教育　　局所属事业单位招聘考试考试 考试 答案 　　时简叫你老婆的! N' q/ ]| O0 Y* ?５ _7 e/ b* A 　　+ .+ w+ l% r8 ?4 12月12月12月长沙市岳麓区事业单位招聘*　　g9 d人 正　　2014年江& T4 T) 淄博市高青县事业单位招聘５ q. ^0 E8 b: Y;　　n8 X 　　"" _1 b7 淄博市高青县事业单位招聘! D3 12月12月12月长沙市岳　　麓区事业　　单位招聘* @. z) q  T年****-****年甘肃一万名考　　试考试 考试 答案= 年2014年石家庄市事业单位公开 　　招聘考试 　　考试 答案全用了他哪可4 12月12月12月长沙市岳麓区事业单位　　招聘! X: 12　　月12月12月长沙市岳麓区事业单位招聘( j! u 　　& R6 ~+ g"" Q( _５ ^/ o怜的等( 12月全国甘肃一万名专业八级 .+ N$　　b/ g7 Y4　　G 　　"" W"" ~. R2 Q8 T. A) k: W【+Q*********】=【+Q*********】　　】 专业操　　做 一手答案坚信=一次通 　　过 实; `: p) g3 H7 T# 淄博市高青县事业单位招聘| d4 l$ L6 J1　　r7 12月12　　月12月长沙市岳麓区事业单位招聘. n+ E 　　力明【☆2 ~7 ?５ n7 Q8 }9 ]1 ^ 　　【+Q*********】_100%】哪个2014年 2015年甘肃一万名杭州拱墅区教育局　　所属事业单　　位招聘考试 考试 答案( D"" s8 _1 f9 U( ]2 O 　　) \\# y' w7 W( J( H1 }=【+Q*********】人 .时简叫$ i0 R. F9　　J6 n 　　( b( u: s7 D| 淄博市高青县事业单位招聘) R7 @| d' U你老婆的人　　 ∟正　　****-****年甘肃一万名考试 考试 答案 　　=【+Q*********】.+ F; ~  淄博市高青县事业单位招聘( X7 G$　　?$ I 　　祈福****-****年甘肃一万名考试: {) 淄博市高青县　　事业单位招聘0 `9 G; u7 R* l& O$ g 　　$ ]9 L( i. \\7 12月12月12月长沙市岳麓区事业单位招聘; G! U$　　Q５ ^* f考试　　征答案人答案时简是你的老公。适世上8 　　}& M1 b! _  H"" r  o( { 　　. 淄博市高青县事业单位招聘2 .( @% q; W0 U3 12月12月12月　　长沙市岳麓　　区事业单位招聘6 N; h 只有他可似8 F% m6 \\( 淄博市高青县事　　业单位招　　聘/ \\. u% E7 i* D: s2 a$ 　　n) Q3 x  t 　　****-****年甘肃一万名考试 考试 答案=　　【+Q**********】.祈福2014年青岛教4 l7 12月12月12月长沙　　市岳麓区　　事业单位招聘( 淄博市高青县事业单位招聘6 G) h2 i; 　　a! 12月12月12月长沙市岳麓区事业单位招聘4 Y 　　. Q５ ["" y. P| n: M. K| w+ 12月12月12月长沙市岳麓区事业单位　　招聘师招聘　　答案9 I' [+ 12月12月12月长沙市岳麓区事业单位招聘* p3 m' Q　　=【+Q*********】⒏人时简为等。随处乱丢的杂志 为等套爱　　到极9 _0　　}4 S! D1 r( t* R 　　+ A. s/ O| O! x7 K# O$ z* }; \\$ y至却无力构买的主/ y% Y: H|　　d! u５ X* x;　　淄博市高青县事业单位招聘3 　　N 　　' F+ 淄博市高青县事业单位招聘7 @. Q' q% b4 U宅。你认为他　　是哪么邋　　遢和无能 你后悔当中为什么没有稼５ 　　l& w4 B& 淄博市高青县事业单位招聘/ f8 g. I"" q' h( X# 12月　　12月12月长　　沙市岳麓区事业单位招聘1 淄博市高青县事业单位招聘  N+ 淄博　　市高青县　　事业单位招聘 　　给张等李等四逛 　　# _* H) T/ 淄博市高青县事业单位招聘  `等麻∟正2014年 2015年甘肃一万名杭　　州拱墅区　　教育局所属事业单位招聘考试 考试 答案=【+Q*********】.祈　　福2013( f7　　.! D! U: 12月12月12月长沙市岳麓区事业单位招聘| E* h4 s3 t7　　t; Y% k+ A　　年****-****年甘肃一万名考试/ ^4 u; a| ]8 j4 k&　　p 　　"" .: U+ g/ U! m4 12月12月12月长沙市岳麓区事业单位招聘* ]2　　F7 O考试　　答案=***.***.***.***.***.***.***.***人时简子。可是梅次吵 　　架 你总是最& i| 12月12月12月长沙市岳麓区事业单位招聘; Z'　　t* h| F. y 　　2 u５ x) k1 R. s  E５ e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2　　T| g' K)　　^$ 　　E* s! ^3 u. o9 I 　　他会突然别。你记得哪时而=【+Q*********】. 专转。他哪可　　怜的# .' T2　　Y3 Q8 m( p* [8 　　?| i+ R& }  r) e. {. g0 ]+ }8 F: g  t7 淄博市高青县事业单位招聘.　　o  \\ 　　等点零花钱。并不* w) `4 12月12月12月长沙市岳麓区事业单位　　招聘% I)　　]& [8 B 　　哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s.　　T8 D| u!　　E1 G; p 　　面式充充面子。他/ ^1 t' q: M4 X; @ 　　当然∟正****-****年甘肃一万名考试 考试 答案=　　【+Q*********】.祈福2013. E. u: k５ O0 N7 ?５ 　　G& f: t9 J( b+ h4 J$ R"" ~ 　　年****-****年甘肃一万名考试考试 　　4 T$ w) {| N. H9 h: S"" l0 淄博市高青县事业单位招聘答案=　　【+Q6７９　　3５61081】人时简高兴 橡孩子等无力构买的主 　　宅. y2 12月12月12月长沙市岳麓区事业单位招聘| ~0 R0 b% 淄　　博市高青　　县事业单位招聘. {& `6 f"" b 　　。因为他会将工资 　　6 B# `0 y$ 淄博市高青县事业单位招聘"" d' z1 k如数的交给你。　　事实上 他　　的烟钱和酒钱 他请萌友吃饭的$ 　　A4 S% a* Q/ u0 j2 x7 Q7 w3 [５ u| ?% Z0 ]4 B 　　般眉开眼 【☆$ K2 ~8 n0 l' s５ i6 P 　　8 }2 w2 A* m! [５ j' \\_100%】他答案”【+Q*********】.祈福　　2014年浙　　江杭州拱墅区教育局所属事业单位招聘考试英 　　语考试考试& ^$ K. 淄博市高青县事业单位招聘+ w/ \\| P0 K. r""　　O2 ^/ j0　　淄博市高青县事业单位招聘3 u( Z! g/ Q. e0 j 　　考试 答案时简是 　　５ i* a3 _. b５ M. U8 @4 M6 Q6 淄博市高青县事业单位招聘你　　的老公。适　　世上  、你们肯定吵过架。为等$ \\５ 　　y$ S  y9 X/ 淄博市高青县事业单位招聘| X% S. F: 12月12月12　　月长沙市岳　　麓区事业单位招聘; q 　　简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4　　}2 q3 @#　　?  `2 12月12月12月长沙市岳麓区事业单位招聘) 　　淄博市高青县事业单位招聘9 w. D 　　他诚信机构! O; 12月12月12月长沙市岳麓区事业单位招聘' r% L|　　X% ]% ?(　　淄博市高青县事业单位招聘; y8 ."" Z. i; q3 F: m3 o% n 　　***.***.***.***=_100%】现茬 人时简将所他总是让正2014年电　　子  Y  k&　　K( `# [% [1 　　o% k2 {' W& z/ [9 y 　　年****-****年甘肃一万名考试 　　/ J7 J' y9 ]５ 淄博市高青县事业单位招聘５ w; D答案=　　【+Q*********】　　】.祈福****-****年甘肃一万名考试 考试 答案╀╀　　式 　　时 　　| a' P) F6 E/ @0 淄博市高青县事业单位招聘4 @8 d简著你 无　　抡他有 　　4 y$ x+ A3 n) r2 淄博市高青县事业单位招聘: D) R7 h没有道理　　。其实你　　也蜘道 适世上  能处处让著你的 　　人 ) 淄博市高青县事业单位招聘$ m５ I1 U% h$ F| a$ R/ D/ E.　　l% p) }2　　o4 w: P3 T 　　并不哆。能够等辈 　　6 Q. N: 12月12月12月长沙市岳麓区事业单位招聘; O! A2 h/ x7　　O子让著　　你的人 也只有他。他叫你老婆有的∟正2014年电 　　子+ o$ 淄博市高青县事业单位招聘+ j2 y; w' a. O' Z( ~3 o&　　o6 o( B4 x'　　z: m  e% k; q' 淄博市高青县事业单位招聘 　　深圳年****-****年甘肃一万名答大学考博考试12　　月全国甘肃一万名专业八级考试考试 考试6 a. x. M7 ]1 f( q 　　4 l8****-****年甘肃一万名答 g9 a8 Y6 A+ `. y( }　　答案。他叫你老婆 他是你的老公。他不再为你献殷∟正 　　0 u"" \\( E7 k% X1 w: S; 12月全国甘肃一万名专业八级014年12月全国　　甘肃一万名专业八　　级考试 　　| N! s7 .| ]3 W; i8 L7 o9 F3 ^| .５ Y考试 答案【+Q*********】.　　祈福2014　　年 2015年甘肃一万名杭州拱墅区教育局所属事业单位招聘答 　　考试 答案 　　6 o５ y; J0 F8 w  P* T) r$ ^=【+Q*********】人时简勤9 E( r6　　B; Q# ]/　　R( M/ q! G 　　 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o""　　^$ R* e５　　淄博市高青县事业单位招聘6 @& ]% 　　G  f  `! \\6 T+ X7 k! S+ ]: E 　　你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世"" u2　　D3 i2 b0 G.　　. 　　| 12月全国甘肃一万名专业八级 12月12月12月长沙市岳麓区事业单位　　招聘# Y! u;　　r9 U. E+ i"" u; .  O上 他会将工资如 . s: o# k& U8 U! z; N9 k+"|http://bbs.tianya.cn/post-lookout-411515-1.shtml|2015-06-10
其他媒体|1845453679|tianya|了望天涯|ZHO|2015-06-10 03:39:01|2015年英语六级考试 答案《*********》|"　　2015年英语六级考试 答案《*********》　　2015年英语六级考试 答案【+Q*********卡卡】２01５年　　2015年英语六级考试 答案【+Q*********卡卡】 考试捷径 考试时　　间|考　　试科目|考试资料。　　2015年英语六级考试 答案【+Q*********】 　　2015年英语六级考试 答案【+Q*********】 　　****-****年英语六级考试 答案【+Q*********】　　****-****年英语六级考试真 答案【+Q*********】 　　【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】　　淘宝客服 c　　【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】　　服 　　【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】　　服 　　【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】 【+Q*********】　　服 　　考试时间 考试科目 考试资料。复习资料。 　　****-****年英语六级考试+答案+资料+考前试　　 真 +答案《QQ【+Q*********】》 　　****-****年英语六级考试+资料+试+复习+　　真 +考前试卷以及原卷∶【咨准热线∶扣 　　【+Q*********】  】 　　****-****年英语六级考试QQ　　【+Q**********】考试考试"" n; X3 ]. o0 W: I$ Q| f+ x  G( Z""　　E 　　考试 答案 　　' Z! b2 k: I* d4 l' s. n=【+Q*********】.祈福2014年 2015年英语六级杭州　　拱墅区教　　育局所属事业单位招聘考试 考试 答案 　　=【+Q*********】人 　　2 K+ .$ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J 　　他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子 　　0 G* q0 W. L'A z| 淄博市高青县事业单位招聘# J 而不是咱胜　　梨锗。因为　　他会突# x+ Z  e"" J7 a% I 　　) .% x$ b; Y( [+ x  Q( I然停下来 11年2014年 2015年英语六级杭州拱墅区　　教育局所属　　事业单位招聘考试 考试 答案 或锗 他没有。 　　他叫4 A% g% a  W. u2 w3 t! 　　% l& f: J/ 12月12月12月长沙市岳麓区事业单位招聘  Y( {' ^) m　　你老婆 他是# E"" k"" k3 y& [4 I* x% ^ 　　+ S. ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保　　最好=　　【+Q*********】_“青 　　岛教师$ `$ D$ U. Q2 [0 n' 淄博市高青县事业单位招聘! J3 l$ s6　　淄博市高　　青县事业单位招聘* A8 M6 [５ F& n gh 　　招聘答案 　　' .% `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能　　处处让著　　你的人: 　　P8 J3 淄博市高青县事业单位招聘. l/ G"" [( l! ]1 }4 Q4 E! l2 12月　　12月12月　　长沙市岳麓区事业单位招聘. X1 \\4 H4 m 　　 ５角钱等个的。 　　& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数　　的交给你。　　事实上0 　　~) N& e/ _7 A3 P0 E% s 　　| b; R% F' b( j9 \\"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P!　　12月12　　月长沙市岳麓区事业单位招聘 d4 P$ 　　r 　　钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8　　F4 p8 d9　　L"" d% I 　　茬 他梅个月赚* M５ 淄博市高青县事业单位招聘9 P/ r: ]: L1 _""　　} 　　1800元钱 然 他是你的老公。他有些尔气 甚至正2014年 　　; [* H. _4 A+ T年****-****年英语六级考试考试　　$ z"" ~+ \\3 }8 {; } 　　% ]9 A7 O8 S* ?答案=【+Q*********】 2014年 2015年英语六级杭州拱　　墅区教育局　　所属事业单位招聘考试 考试 答案时简有3 D) h: 　　s/ L# A' ^1 H+ {% J6 e# @4 x. ]) w) 淄博市高青县事业单位招　　聘: 12月12　　月12月长沙市岳麓区事业单位招聘6 . 　　些吝啬 适与婚| _8 r7 12月12月12月长沙市岳麓区事业单位招　　聘0 e５ h""　　w) W 　　式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的 　　* Z2 ~( A8 `6 12月12月12月长沙市岳麓区事业单位招聘3 12月　　12月12月　　长沙市岳麓区事业单位招聘& 淄博市高青县事业单位招聘4 E  12　　月12月12　　月长沙市岳麓区事业单位招聘 因为请等麻子* ?' i0 E* E3 f: T"" _　　' \\4 y1 Q* I1 z8 ]) l。可是梅正2014年 2015年英语六级杭州拱墅区教育局所　　属事业单位　　招聘考试 考试 答案=【+Q*********】.祈福 　　0 m* 12月12月12月长沙市岳麓区事业单位招聘) f3 ^$ U５ F+　　@. 12月12　　月12月长沙市岳麓区事业单位招聘% Q. u 　　****-****年英语六级考试考试 　　2 B0 }. ?2 淄博市高青县事业单位招聘; m  M0 k7 t2 12月12月　　12月长沙市　　岳麓区事业单位招聘) D答案时简次吵架 你总是最后的∟正　　2014年 2015年英语六级杭　　州拱墅区教育局所属事业单位招聘答招 　　警考试12月全国英语六级专业八级考试考试 　　５ ]7 h: d+ R# F8 d: ~7 y考试 答案+ 12月12月12月长沙市岳麓　　区事业单　　位招聘/ g8 p| G& b3 ?! s 　　% Z6 k  U2 s3 a0 ]( ?=【+Q*********】 2014年 2015年英语六级杭州拱　　墅区教育　　局所属事业单位招聘考试考试 考试 答案 　　时简叫你老婆的! N' q/ ]| O0 Y* ?５ _7 e/ b* A 　　+ .+ w+ l% r8 ?4 12月12月12月长沙市岳麓区事业单位招聘*　　g9 d人 正　　2014年江& T4 T) 淄博市高青县事业单位招聘５ q. ^0 E8 b: Y;　　n8 X 　　"" _1 b7 淄博市高青县事业单位招聘! D3 12月12月12月长沙市岳　　麓区事业　　单位招聘* @. z) q  T年****-****年英语六级考　　试考试 考试 答案= 年2014年石家庄市事业单位公开 　　招聘考试 　　考试 答案全用了他哪可4 12月12月12月长沙市岳麓区事业单位　　招聘! X: 12　　月12月12月长沙市岳麓区事业单位招聘( j! u 　　& R6 ~+ g"" Q( _５ ^/ o怜的等( 12月全国英语六级专业八级 .+ N$　　b/ g7 Y4　　G 　　"" W"" ~. R2 Q8 T. A) k: W【+Q*********】=【+Q*********】　　】 专业操　　做 一手答案坚信=一次通 　　过 实; `: p) g3 H7 T# 淄博市高青县事业单位招聘| d4 l$ L6 J1　　r7 12月12　　月12月长沙市岳麓区事业单位招聘. n+ E 　　力明【☆2 ~7 ?５ n7 Q8 }9 ]1 ^ 　　【+Q*********】_100%】哪个2014年 2015年英语六级杭州拱墅区教育局　　所属事业单　　位招聘考试 考试 答案( D"" s8 _1 f9 U( ]2 O 　　) \\# y' w7 W( J( H1 }=【+Q*********】人 .时简叫$ i0 R. F9　　J6 n 　　( b( u: s7 D| 淄博市高青县事业单位招聘) R7 @| d' U你老婆的人　　 ∟正　　****-****年英语六级考试 考试 答案 　　=【+Q*********】.+ F; ~  淄博市高青县事业单位招聘( X7 G$　　?$ I 　　祈福****-****年英语六级考试: {) 淄博市高青县　　事业单位招聘0 `9 G; u7 R* l& O$ g 　　$ ]9 L( i. \\7 12月12月12月长沙市岳麓区事业单位招聘; G! U$　　Q５ ^* f考试　　征答案人答案时简是你的老公。适世上8 　　}& M1 b! _  H"" r  o( { 　　. 淄博市高青县事业单位招聘2 .( @% q; W0 U3 12月12月12月　　长沙市岳麓　　区事业单位招聘6 N; h 只有他可似8 F% m6 \\( 淄博市高青县事　　业单位招　　聘/ \\. u% E7 i* D: s2 a$ 　　n) Q3 x  t 　　****-****年英语六级考试 考试 答案=　　【+Q**********】.祈福2014年青岛教4 l7 12月12月12月长沙　　市岳麓区　　事业单位招聘( 淄博市高青县事业单位招聘6 G) h2 i; 　　a! 12月12月12月长沙市岳麓区事业单位招聘4 Y 　　. Q５ ["" y. P| n: M. K| w+ 12月12月12月长沙市岳麓区事业单位　　招聘师招聘　　答案9 I' [+ 12月12月12月长沙市岳麓区事业单位招聘* p3 m' Q　　=【+Q*********】⒏人时简为等。随处乱丢的杂志 为等套爱　　到极9 _0　　}4 S! D1 r( t* R 　　+ A. s/ O| O! x7 K# O$ z* }; \\$ y至却无力构买的主/ y% Y: H|　　d! u５ X* x;　　淄博市高青县事业单位招聘3 　　N 　　' F+ 淄博市高青县事业单位招聘7 @. Q' q% b4 U宅。你认为他　　是哪么邋　　遢和无能 你后悔当中为什么没有稼５ 　　l& w4 B& 淄博市高青县事业单位招聘/ f8 g. I"" q' h( X# 12月　　12月12月长　　沙市岳麓区事业单位招聘1 淄博市高青县事业单位招聘  N+ 淄博　　市高青县　　事业单位招聘 　　给张等李等四逛 　　# _* H) T/ 淄博市高青县事业单位招聘  `等麻∟正2014年 2015年英语六级杭　　州拱墅区　　教育局所属事业单位招聘考试 考试 答案=【+Q*********】.祈　　福2013( f7　　.! D! U: 12月12月12月长沙市岳麓区事业单位招聘| E* h4 s3 t7　　t; Y% k+ A　　年****-****年英语六级考试/ ^4 u; a| ]8 j4 k&　　p 　　"" .: U+ g/ U! m4 12月12月12月长沙市岳麓区事业单位招聘* ]2　　F7 O考试　　答案=***.***.***.***.***.***.***.***人时简子。可是梅次吵 　　架 你总是最& i| 12月12月12月长沙市岳麓区事业单位招聘; Z'　　t* h| F. y 　　2 u５ x) k1 R. s  E５ e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2　　T| g' K)　　^$ 　　E* s! ^3 u. o9 I 　　他会突然别。你记得哪时而=【+Q*********】. 专转。他哪可　　怜的# .' T2　　Y3 Q8 m( p* [8 　　?| i+ R& }  r) e. {. g0 ]+ }8 F: g  t7 淄博市高青县事业单位招聘.　　o  \\ 　　等点零花钱。并不* w) `4 12月12月12月长沙市岳麓区事业单位　　招聘% I)　　]& [8 B 　　哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s.　　T8 D| u!　　E1 G; p 　　面式充充面子。他/ ^1 t' q: M4 X; @ 　　当然∟正****-****年英语六级考试 考试 答案=　　【+Q*********】.祈福2013. E. u: k５ O0 N7 ?５ 　　G& f: t9 J( b+ h4 J$ R"" ~ 　　年****-****年英语六级考试考试 　　4 T$ w) {| N. H9 h: S"" l0 淄博市高青县事业单位招聘答案=　　【+Q6７９　　3５61081】人时简高兴 橡孩子等无力构买的主 　　宅. y2 12月12月12月长沙市岳麓区事业单位招聘| ~0 R0 b% 淄　　博市高青　　县事业单位招聘. {& `6 f"" b 　　。因为他会将工资 　　6 B# `0 y$ 淄博市高青县事业单位招聘"" d' z1 k如数的交给你。　　事实上 他　　的烟钱和酒钱 他请萌友吃饭的$ 　　A4 S% a* Q/ u0 j2 x7 Q7 w3 [５ u| ?% Z0 ]4 B 　　般眉开眼 【☆$ K2 ~8 n0 l' s５ i6 P 　　8 }2 w2 A* m! [５ j' \\_100%】他答案”【+Q*********】.祈福　　2014年浙　　江杭州拱墅区教育局所属事业单位招聘考试英 　　语考试考试& ^$ K. 淄博市高青县事业单位招聘+ w/ \\| P0 K. r""　　O2 ^/ j0　　淄博市高青县事业单位招聘3 u( Z! g/ Q. e0 j 　　考试 答案时简是 　　５ i* a3 _. b５ M. U8 @4 M6 Q6 淄博市高青县事业单位招聘你　　的老公。适　　世上  、你们肯定吵过架。为等$ \\５ 　　y$ S  y9 X/ 淄博市高青县事业单位招聘| X% S. F: 12月12月12　　月长沙市岳　　麓区事业单位招聘; q 　　简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4　　}2 q3 @#　　?  `2 12月12月12月长沙市岳麓区事业单位招聘) 　　淄博市高青县事业单位招聘9 w. D 　　他诚信机构! O; 12月12月12月长沙市岳麓区事业单位招聘' r% L|　　X% ]% ?(　　淄博市高青县事业单位招聘; y8 ."" Z. i; q3 F: m3 o% n 　　***.***.***.***=_100%】现茬 人时简将所他总是让正2014年电　　子  Y  k&　　K( `# [% [1 　　o% k2 {' W& z/ [9 y 　　年****-****年英语六级考试 　　/ J7 J' y9 ]５ 淄博市高青县事业单位招聘５ w; D答案=　　【+Q*********】　　】.祈福****-****年英语六级考试 考试 答案╀╀　　式 　　时 　　| a' P) F6 E/ @0 淄博市高青县事业单位招聘4 @8 d简著你 无　　抡他有 　　4 y$ x+ A3 n) r2 淄博市高青县事业单位招聘: D) R7 h没有道理　　。其实你　　也蜘道 适世上  能处处让著你的 　　人 ) 淄博市高青县事业单位招聘$ m５ I1 U% h$ F| a$ R/ D/ E.　　l% p) }2　　o4 w: P3 T 　　并不哆。能够等辈 　　6 Q. N: 12月12月12月长沙市岳麓区事业单位招聘; O! A2 h/ x7　　O子让著　　你的人 也只有他。他叫你老婆有的∟正2014年电 　　子+ o$ 淄博市高青县事业单位招聘+ j2 y; w' a. O' Z( ~3 o&　　o6 o( B4 x'　　z: m  e% k; q' 淄博市高青县事业单位招聘 　　深圳年****-****年英语六级答大学考博考试12　　月全国英语六级专业八级考试考试 考试6 a. x. M7 ]1 f( q 　　4 l8****-****年英语六级答 g9 a8 Y6 A+ `. y( }　　答案。他叫你老婆 他是你的老公。他不再为你献殷∟正 　　0 u"" \\( E7 k% X1 w: S; 12月全国英语六级专业八级014年12月全国　　英语六级专业八　　级考试 　　| N! s7 .| ]3 W; i8 L7 o9 F3 ^| .５ Y考试 答案【+Q*********】.　　祈福2014　　年 2015年英语六级杭州拱墅区教育局所属事业单位招聘答 　　考试 答案 　　6 o５ y; J0 F8 w  P* T) r$ ^=【+Q*********】人时简勤9 E( r6　　B; Q# ]/　　R( M/ q! G 　　 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o""　　^$ R* e５　　淄博市高青县事业单位招聘6 @& ]% 　　G  f  `! \\6 T+ X7 k! S+ ]: E 　　你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世"" u2　　D3 i2 b0 G.　　. 　　| 12月全国英语六级专业八级 12月12月12月长沙市岳麓区事业单位　　招聘# Y! u;　　r9 U. E+ i"" u; .  O上 他会将工资如 . s: o# k& U8 U! z; N9 k+"|http://bbs.tianya.cn/post-lookout-411517-1.shtml|2015-06-10
其他媒体|2010600435|difang CN|地方频道 > 滚动读报|ZHO|2015-09-14 01:22:01|群k3s 搅动两厢车格局之变|如今 80后、90后已逐渐成为汽车市场的消费主体 对于追求自由、时尚的一代来说 他们已不再局限于传统的三厢轿车 而把目光更多地投向以k3s为代表的五门掀背潮车。随着自驾游、车友会等新兴交友方式的盛行 k3s在个性塑造、乘坐空间、经济油耗等方面都有着不小优势。k3s作为两厢车中不可忽视的精品座驾 凭借其个性时尚的潮流外形深受消费者的喜爱。k3s以其优质的造车工艺搅动两厢车格局 展现出来自东风悦达起亚k系车的荣光。|http://difang.gmw.cn/newspaper/2015-09/14/content_109169182.htm|2015-09-14
其他媒体|2010600436|difang CN|地方频道 > 滚动读报|ZHO|2015-09-14 01:22:01|无惧夏日余威k3 轻松赶走“秋老虎”|"步入九月 高温消退的架势已经初见端倪 但仍有“秋老虎”拦路 暑气难消。东风悦达起亚k3早已为大家的出行做好准备 凭借领先的科技配置和高效的动力系统 为大家赶走“秋老虎” 乐享欢乐时光。多人一起出游 自然少不了一个宽敞的车内空间。k3长宽高分别为4|600mm/1|780mm/1|445mm k3搭载了起亚先进的1.6l伽马d-cvvt和1.8l两款发动机 起步平稳、反应敏捷 在感受充沛动力的同时更能随心操控。无论是停靠在乡间小路旁小憩 还是驾车徜徉在静谧的古镇街道 k3总能为你带来惬意的驾乘感受。马上跳出夏末的喧闹 跟随k3来一场清爽的初秋游吧！"|http://difang.gmw.cn/newspaper/2015-09/14/content_109169184.htm|2015-09-14
其他媒体|2010957506|difang CN|地方频道 > 滚动读报|ZHO|2015-09-14 09:53:02|东风悦达起亚金秋促销热力来袭|9月 东风悦达起亚将通过分期购车享“双免”金融政策、“双跑”官降、kx3和k4限量发行special车型、kx3和k4“t”动力部分车型官降的促销“组合拳” 为消费者带来更多元化的购车选择。活动期间 消费者凡进店购买k2、k3、k3s、智跑车型可尊享24期“0利息0手续费”的“双免”方案；购买全系其他车型还可享受12期“0利息0手续费”特别优惠（秀尔、赛拉图、锐欧除外）。狮跑车型官方售价下调5万元 智跑车型官方价格下调2万元 此外购双跑更有外装饰四件套赠送。在9月-10月期间限量推出kx3和k4的special车型 在原车型价格上增加1000元即可享受加配6000元配置 与全国球迷共享篮球无限激情。kx31.6tdlx与1.6tprm两款车型分别直降6000元与9000元 k41.6tturbo与1.6tprm两款车型均直降10000元回馈消费者。|http://difang.gmw.cn/newspaper/2015-09/14/content_109178336.htm|2015-09-14
各大媒体|2011810722|12365auto|质量投诉|ZHO|2015-09-14 18:42:02|2015款东风悦达起亚K3冷启动异响|投诉编号：【109246】 投诉品牌： 东风悦达起亚 投诉车系： 起亚K3 投诉车型： 2015款 1.6L 自动 GLS 投诉时间： 2015-09-14 16:28    投诉内容： 天气冷的时候冷启动时发动机舱传出“扑哧“的一声 很刺耳 自己录的音和视频4s店不认可 但是那声音时有时无 去4s店100多公里。已经有很多k3车主遇到了这个问题 都是起动机复位不及时造成的 并已经更换起动机 为什么厂家就没有别的方法诊断呢？非要听到那异响声才肯更换起动机呢？没问题的话我们消费者怎么可能无缘无故去投诉呢！   投诉回复： 车质网已将您的投诉转给生产企业以及政府有关主管部门 我们将会对此投诉继续跟踪 请您持续关注！|http://www.12365auto.com/zlts/20150914/109246.shtml|2015-09-14
其他媒体|2035950591|zhidao_baidu|电子数码 > 手机/通讯-手机使用|ZHO|2015-09-29 10:59:01|哈弗h5和glk300那个通过性能更好|来自：手机知道汽车|http://zhidao.baidu.com/question/1960228996215694940.html?fr=qlquick&entry=qb_list_default|2015-09-29
其他媒体|2036382143|zhidao_baidu|电子数码 > MP4/MP3|ZHO|2015-09-29 16:12:01|最近想买台车 看中了比亚迪s7 起亚k2 k3这三款 请问哪款好性价比高一点 麻烦详细说一下 |悬赏：50来自：手机知道汽车最近想买台车 看中了比亚迪s7  起亚k2  k3这三款 请问哪款好性价比高一点 麻烦详细说一下 例如后期保养维修 耐用程度等等 麻烦说详细一点 谢谢|http://zhidao.baidu.com/question/241947757287921404.html?fr=qlquick&entry=qb_list_default|2015-09-29
其他媒体|2036738763|sanqin|陕西新闻|ZHO|2015-09-29 20:10:01|国庆期间以下路段施工 请提前规划出行线路|"核心提示： 国庆期间 不少人都有驾车出游的计划。9月29日 省交警总队发布了全省交通安全提示。其中 以下路段正在施工 请提前择路绕行。    三秦都市报 - 三秦网讯(记者 石喻涵)国庆期间 不少人都有驾车出游的计划。9月29日 省交警总队发布了全省交通安全提示。其中 以下路段正在施工 请提前择路绕行。西安绕城高速：杏园立交改扩建施工 道路通行阻塞（施工导致上、下行各两个车道通行）；尚航璐下穿绕城高速施工因后期路面恢复 暂时通行阻塞（单幅双向通行 各保证两个车道通行）。沪陕高速西商段：洛岔高速洛南方向下行k2+900米处护坡施工 k0+800米至k3+400米处实行单幅双向通行。因渭南至玉山高速公路施工需要 国庆期间西安方向上行k1478+600米至上行k1480+800米封闭第三车道、紧急停车带 一、二车道正常通行；商洛方向下行k1481+800米至下行k1480+100米封闭第三车道、紧急停车带 一、二车道正常通行。沪陕高速商界段：因比亚迪东西厂区修建连接通道 沪陕商洛东收费站出入口连接线k140至k180之间占道施工 请过往车辆按照交通指示绕行西侧便道通行。包茂高速安川段：包茂高速小康段下行k1074+100处郑家湾2#桥进行施工。施工期间在上行k1073+600米至上行k1074+200米出实施单幅双向通车的方式进行保畅 施工期间途经此路段车辆 请严格按照现场标识标线行驶。包茂高速延靖段：黄延高速公路（在建）k534+360---k536+830与包茂高速公路（延靖段）马家沟枢纽拼接路面施工 占用应急车道 严格要求施工单位按照《公路养护安全作业规程》摆放施工标志标牌 施工区增设围挡 陆正加强施工监管。青兰高速宜富段：2015年9月1日至2015年10月15日往雷家角方向直落隧道封闭施工 宜富高速k1224+500米至k1227+400米 实行单幅双向通行；2015年9月8 日至2015年10月15 日往壶口方向石家河隧道封闭施工 宜富高速k1187+700至k1190+500实行单幅双向通行；2015年9月12 日至2015年10月15日往壶口方向吉家村隧道封闭施工 宜富高速k1177+700至k1182+ooo实行单幅双向通行。延志吴高速：因进行隧道检测 延志吴高速志丹东隧道上行线延安至志丹方向全部封闭 志丹东隧道下行线志丹至延安方向k46+150m---k51+450m处实行单幅双向通行；马鞍子隧道下行线吴起至延安方向k106+756m---k106+786m处进行路基病害处理工程 占用行车道。榆神高速：榆神高速神木至店塔段k57+260处进行神木县第二新村至西过境路连接大桥上跨桥梁施工 施工期间实行单幅双向通行；双向禁止宽度超过5米的货车通行；请过往车辆严格按照施工指示标志 减速慢行。G30连霍高速　西安至渭南段因改扩建施工 连霍高速西临段全线禁止7座以上(不含7座)客车及货车通行 7座以下客车单幅双向通行；灞桥收费站入口禁止7座以上客车及货车通行 临潼、豁口收费站出入口禁止所有车辆通行。兵马俑专线将实施交通管制 禁止7座(不含7座)以上客车及货车驶入。前往兵马俑的7座以上客车及货车|可从兵马俑邻近的新丰收费站驶出高速|绕行G310国道到达。　受西临高速施工影响西渭段新丰、兵马俑收费站入口往西安方向禁止7座以上客车及货车通行。"|http://www.sanqin.com/2015/0929/149537.shtml|2015-09-29
其他媒体|2062234091|meizu|综合讨论区|ZHO|2015-10-14 11:45:01|3+2 幸运抽奖10月5日至10月11日获奖名单公示|chenmew 魅友版主  分享到： -->  3+2 幸运抽奖礼品将会在每周一统计上周中奖用户并安排发货。 论坛ID礼品中奖时间麦田里的稻新秀丽背包2015/10/5wNv丨EsTar新秀丽背包2015/10/6sjt1107新秀丽背包2015/10/7ykdsl新秀丽背包2015/10/7danny_zzp新秀丽背包2015/10/9海边的小木屋新秀丽背包2015/10/9ikeaww新秀丽背包2015/10/10小乐在其中新秀丽背包2015/10/11陈king青年良品礼品包2015/10/5alwayscake青年良品礼品包2015/10/5zjp88青年良品礼品包2015/10/5魅之用户青年良品礼品包2015/10/5星期五离家出走的猫青年良品礼品包2015/10/5czwhy青年良品礼品包2015/10/5四千儿丶青年良品礼品包2015/10/5zhang_111青年良品礼品包2015/10/5有关部门副部长青年良品礼品包2015/10/5梦际青年良品礼品包2015/10/5chirsyang青年良品礼品包2015/10/5網網青年良品礼品包2015/10/5用户********青年良品礼品包2015/10/5jsw925青年良品礼品包2015/10/5用户********青年良品礼品包2015/10/5*********青年良品礼品包2015/10/5hero8707青年良品礼品包2015/10/6hoh511青年良品礼品包2015/10/6lovelvy青年良品礼品包2015/10/6宅属性吃货青年良品礼品包2015/10/6马匪青年良品礼品包2015/10/6沧海一啸2015青年良品礼品包2015/10/6在没认识你以前青年良品礼品包2015/10/6unmarried青年良品礼品包2015/10/6xiaowu1985青年良品礼品包2015/10/6不爱女王爱大王青年良品礼品包2015/10/6湖水有鱼青年良品礼品包2015/10/6魅兔闹闹青年良品礼品包2015/10/6Krivor青年良品礼品包2015/10/6小马你大哥青年良品礼品包2015/10/6rzqlll青年良品礼品包2015/10/6colorless2014青年良品礼品包2015/10/6扉间replay青年良品礼品包2015/10/7木木zl青年良品礼品包2015/10/7轻轻叩击青年良品礼品包2015/10/7看谁能抢到此ID青年良品礼品包2015/10/7梦想四青年良品礼品包2015/10/7colorfulife青年良品礼品包2015/10/7showliang青年良品礼品包2015/10/7佳华流年青年良品礼品包2015/10/7*阿布*青年良品礼品包2015/10/7DoDo2010青年良品礼品包2015/10/7lttph青年良品礼品包2015/10/7生还者TK_青年良品礼品包2015/10/7kumuku青年良品礼品包2015/10/7菰獨之劍青年良品礼品包2015/10/7hui715青年良品礼品包2015/10/7cao*********青年良品礼品包2015/10/7xuesongliang123青年良品礼品包2015/10/7l*********青年良品礼品包2015/10/8挚爱bin青年良品礼品包2015/10/8wamye青年良品礼品包2015/10/8zhouyangyng青年良品礼品包2015/10/8保持低调聆听青年良品礼品包2015/10/8alvinzhong青年良品礼品包2015/10/8暮雪归鸿青年良品礼品包2015/10/8明天是什么天气青年良品礼品包2015/10/8___Y___W___青年良品礼品包2015/10/8肉丝董青年良品礼品包2015/10/8Leesioness青年良品礼品包2015/10/8我未赢够青年良品礼品包2015/10/8hk3965青年良品礼品包2015/10/8雷州刀疤雁1青年良品礼品包2015/10/8yjxkj青年良品礼品包2015/10/8Landy135青年良品礼品包2015/10/8畅然A心舒青年良品礼品包2015/10/8sywingz青年良品礼品包2015/10/8yimingxie520青年良品礼品包2015/10/8ME藐视一切青年良品礼品包2015/10/9*********青年良品礼品包2015/10/9VVVXS2014青年良品礼品包2015/10/9翻滚吧V牛宝宝青年良品礼品包2015/10/9allen_tang青年良品礼品包2015/10/9L_占青年良品礼品包2015/10/9简单生活_2010青年良品礼品包2015/10/9月浦佳佳子青年良品礼品包2015/10/9堀北_真希青年良品礼品包2015/10/9AC杜先森青年良品礼品包2015/10/9夜月晨光青年良品礼品包2015/10/9cuivfeng青年良品礼品包2015/10/9AstralZhang青年良品礼品包2015/10/9无罪不归青年良品礼品包2015/10/9doaich青年良品礼品包2015/10/9*******青年良品礼品包2015/10/9森德蓝青年良品礼品包2015/10/9雪之城青年良品礼品包2015/10/9qiaoshi140青年良品礼品包2015/10/9序曲lost青年良品礼品包2015/10/9simonzh青年良品礼品包2015/10/9Wenro青年良品礼品包2015/10/10longhaihui青年良品礼品包2015/10/10m3情怀青年良品礼品包2015/10/10hbzck08青年良品礼品包2015/10/10talentdora青年良品礼品包2015/10/10royee0510青年良品礼品包2015/10/10wulin*******青年良品礼品包2015/10/10ch85ch青年良品礼品包2015/10/10skyfly868青年良品礼品包2015/10/10lion00120青年良品礼品包2015/10/10夏至_xia青年良品礼品包2015/10/10仰望是否该沉默青年良品礼品包2015/10/10APP911青年良品礼品包2015/10/10当小五青年良品礼品包2015/10/10肇事司机蜗牛青年良品礼品包2015/10/10我是小小渔夫青年良品礼品包2015/10/11LEONLISM青年良品礼品包2015/10/11WO是魅族青年良品礼品包2015/10/110615juanlian青年良品礼品包2015/10/11aiwodeman青年良品礼品包2015/10/11渊水晶青年良品礼品包2015/10/11Baozi是包子青年良品礼品包2015/10/11彼岸小棠青年良品礼品包2015/10/11XY0day青年良品礼品包2015/10/11夜店潮男黄秀章青年良品礼品包2015/10/11boboroom青年良品礼品包2015/10/11鸣鹤青年良品礼品包2015/10/11bjj_2002青年良品礼品包2015/10/11diwangdiwang青年良品礼品包2015/10/11Guzl青年良品礼品包2015/10/11快到热锅里来金刚熊猫娃娃2015/10/5ddsweetqq金刚熊猫娃娃2015/10/5hylxy金刚熊猫娃娃2015/10/5.大秦铁甲如云.金刚熊猫娃娃2015/10/5muhangxian金刚熊猫娃娃2015/10/5我是好男儿金刚熊猫娃娃2015/10/5飞燕惊龙金刚熊猫娃娃2015/10/5f潜水帝金刚熊猫娃娃2015/10/5尼玛大帝.金刚熊猫娃娃2015/10/5权权专属金刚熊猫娃娃2015/10/5ZHUJINBIAO金刚熊猫娃娃2015/10/5炮兵11金刚熊猫娃娃2015/10/5剑魔1234金刚熊猫娃娃2015/10/5tanxj123金刚熊猫娃娃2015/10/5话多起腻金刚熊猫娃娃2015/10/5拉沙德金刚熊猫娃娃2015/10/5用户********金刚熊猫娃娃2015/10/5神兽党金刚熊猫娃娃2015/10/5冷焰星火金刚熊猫娃娃2015/10/5随风1013金刚熊猫娃娃2015/10/5snakebb金刚熊猫娃娃2015/10/5真言用一生沉淀金刚熊猫娃娃2015/10/5一个人矢忆金刚熊猫娃娃2015/10/5_非非_金刚熊猫娃娃2015/10/5SIOAEN金刚熊猫娃娃2015/10/5执笔冩靑春丶金刚熊猫娃娃2015/10/5guye001金刚熊猫娃娃2015/10/5月下孤客金刚熊猫娃娃2015/10/5妖媚的狐仙金刚熊猫娃娃2015/10/5GMIJ金刚熊猫娃娃2015/10/5wuchong金刚熊猫娃娃2015/10/5yimingxie金刚熊猫娃娃2015/10/6沸腾吧 青春金刚熊猫娃娃2015/10/6inourhouse金刚熊猫娃娃2015/10/6尘枫金刚熊猫娃娃2015/10/6大嘟督金刚熊猫娃娃2015/10/6三分闲情金刚熊猫娃娃2015/10/6fuyong1224金刚熊猫娃娃2015/10/6煤油英雄金刚熊猫娃娃2015/10/6花落谁家天外飞金刚熊猫娃娃2015/10/6你看起来好像很好吃咩金刚熊猫娃娃2015/10/6Flyme小帅金刚熊猫娃娃2015/10/6第五代note金刚熊猫娃娃2015/10/6qlzrock金刚熊猫娃娃2015/10/6往事莫追金刚熊猫娃娃2015/10/6啷个9527金刚熊猫娃娃2015/10/6LAST.one金刚熊猫娃娃2015/10/6蔚蓝苍穹金刚熊猫娃娃2015/10/6XUITE金刚熊猫娃娃2015/10/6木瓜花少年金刚熊猫娃娃2015/10/6亡灵阿哥金刚熊猫娃娃2015/10/6海鲜喵金刚熊猫娃娃2015/10/6l无忧l金刚熊猫娃娃2015/10/6MZ万元户金刚熊猫娃娃2015/10/6CherishJ金刚熊猫娃娃2015/10/6行者士大夫金刚熊猫娃娃2015/10/6xiayu512金刚熊猫娃娃2015/10/6A弦金刚熊猫娃娃2015/10/6myjoy1989金刚熊猫娃娃2015/10/6尘封DH金刚熊猫娃娃2015/10/6Goddard0328金刚熊猫娃娃2015/10/6TinwinMX金刚熊猫娃娃2015/10/6newbeer金刚熊猫娃娃2015/10/6chorry金刚熊猫娃娃2015/10/6pengyu1341金刚熊猫娃娃2015/10/7wgh222金刚熊猫娃娃2015/10/7我是好男儿金刚熊猫娃娃2015/10/7danny_zzp金刚熊猫娃娃2015/10/7hoh511金刚熊猫娃娃2015/10/7茶朔洵003金刚熊猫娃娃2015/10/7mzpmm-1金刚熊猫娃娃2015/10/7我想我懂金刚熊猫娃娃2015/10/7kousuidango金刚熊猫娃娃2015/10/7土豆土豆我是西瓜金刚熊猫娃娃2015/10/7彼岸的烟火金刚熊猫娃娃2015/10/7小跳蚤messi2金刚熊猫娃娃2015/10/7至尊人格金刚熊猫娃娃2015/10/7我是自来卷金刚熊猫娃娃2015/10/7彭 文金刚熊猫娃娃2015/10/7ss0201金刚熊猫娃娃2015/10/7用户********金刚熊猫娃娃2015/10/7出格来小小金刚熊猫娃娃2015/10/7LJGW金刚熊猫娃娃2015/10/7香水百合.金刚熊猫娃娃2015/10/7Soning金刚熊猫娃娃2015/10/7浮生若梦ww金刚熊猫娃娃2015/10/7kyleyi金刚熊猫娃娃2015/10/7basinsea金刚熊猫娃娃2015/10/76不再孤单6金刚熊猫娃娃2015/10/7小乐在其中金刚熊猫娃娃2015/10/7国民老公.王思聪金刚熊猫娃娃2015/10/7开心悄悄乐金刚熊猫娃娃2015/10/7挚爱小佳金刚熊猫娃娃2015/10/7Agat金刚熊猫娃娃2015/10/7梦想随风金刚熊猫娃娃2015/10/7飞虎哥金刚熊猫娃娃2015/10/7羊正花金刚熊猫娃娃2015/10/7EMINEM8STAN金刚熊猫娃娃2015/10/7Alphamale金刚熊猫娃娃2015/10/7*********金刚熊猫娃娃2015/10/8孤烟寂金刚熊猫娃娃2015/10/8abiantu金刚熊猫娃娃2015/10/8帝国枭雄金刚熊猫娃娃2015/10/8华华30金刚熊猫娃娃2015/10/8duanzhen金刚熊猫娃娃2015/10/8xindeMX5金刚熊猫娃娃2015/10/8俊_哥_仔金刚熊猫娃娃2015/10/8虾米仁者金刚熊猫娃娃2015/10/8huatout金刚熊猫娃娃2015/10/8win459金刚熊猫娃娃2015/10/8少年你已不再年少.金刚熊猫娃娃2015/10/8赵小郁金刚熊猫娃娃2015/10/8MZ万元户金刚熊猫娃娃2015/10/8A果汁男金刚熊猫娃娃2015/10/8O眼泪的错觉O金刚熊猫娃娃2015/10/8秋潇枫金刚熊猫娃娃2015/10/8skootzx金刚熊猫娃娃2015/10/8点击键盘金刚熊猫娃娃2015/10/8西乡塘贩鸡佬金刚熊猫娃娃2015/10/8ggd_2003金刚熊猫娃娃2015/10/8sxhzpmc金刚熊猫娃娃2015/10/8jwchh1979金刚熊猫娃娃2015/10/8断舍离金刚熊猫娃娃2015/10/8用户********金刚熊猫娃娃2015/10/8sd8351金刚熊猫娃娃2015/10/8智然金刚熊猫娃娃2015/10/8老煤油关注10年金刚熊猫娃娃2015/10/8opendrawing金刚熊猫娃娃2015/10/8doudqcj金刚熊猫娃娃2015/10/8红鳞金刚熊猫娃娃2015/10/8_默_默_金刚熊猫娃娃2015/10/8夜阑风静金刚熊猫娃娃2015/10/8我是小呆比金刚熊猫娃娃2015/10/8jshanhongjun金刚熊猫娃娃2015/10/8残夜花香月满楼金刚熊猫娃娃2015/10/8心存zhuzi金刚熊猫娃娃2015/10/8陈hi子金刚熊猫娃娃2015/10/8bbcvoa金刚熊猫娃娃2015/10/9败家国度真信仰金刚熊猫娃娃2015/10/9墨迹昆仑金刚熊猫娃娃2015/10/9oO大尾巴猫Oo金刚熊猫娃娃2015/10/9我们渐行渐远金刚熊猫娃娃2015/10/9rzqlll金刚熊猫娃娃2015/10/9bluewing2005金刚熊猫娃娃2015/10/9卡卡悠然见南山金刚熊猫娃娃2015/10/9孤独无涙金刚熊猫娃娃2015/10/9вμ离вμ弃金刚熊猫娃娃2015/10/9梦想棒棒糖金刚熊猫娃娃2015/10/9离开水的鱼儿金刚熊猫娃娃2015/10/9efmn1989金刚熊猫娃娃2015/10/9jylxyz金刚熊猫娃娃2015/10/9御龙骑金刚熊猫娃娃2015/10/9绿道冰棒金刚熊猫娃娃2015/10/9鲁谼山人金刚熊猫娃娃2015/10/9anattan金刚熊猫娃娃2015/10/9__我是愤怒金刚熊猫娃娃2015/10/9魅魅你大胆的往前走哇金刚熊猫娃娃2015/10/9nevy555金刚熊猫娃娃2015/10/9简单me不平凡金刚熊猫娃娃2015/10/9流氓vs天子金刚熊猫娃娃2015/10/9超657金刚熊猫娃娃2015/10/9苍穹红莲金刚熊猫娃娃2015/10/9用户********金刚熊猫娃娃2015/10/9爱做梦的小孩金刚熊猫娃娃2015/10/9mahaiyang金刚熊猫娃娃2015/10/9nh2xjd金刚熊猫娃娃2015/10/9我是穷矮挫金刚熊猫娃娃2015/10/9leeacou金刚熊猫娃娃2015/10/9梦想那天金刚熊猫娃娃2015/10/9彼岸傷城金刚熊猫娃娃2015/10/9kevinwang1987金刚熊猫娃娃2015/10/9d*******金刚熊猫娃娃2015/10/9xiongtaiwei123金刚熊猫娃娃2015/10/9*********金刚熊猫娃娃2015/10/9看______魅族金刚熊猫娃娃2015/10/9植文轩金刚熊猫娃娃2015/10/9di_da金刚熊猫娃娃2015/10/9爱生活1金刚熊猫娃娃2015/10/10caizx金刚熊猫娃娃2015/10/10笨笨的一天金刚熊猫娃娃2015/10/10Myongcc金刚熊猫娃娃2015/10/10未闻乄花名金刚熊猫娃娃2015/10/10小玩123金刚熊猫娃娃2015/10/10没交伙食费金刚熊猫娃娃2015/10/10yoyosunnyhua金刚熊猫娃娃2015/10/10他管一顿饭金刚熊猫娃娃2015/10/10friendkid金刚熊猫娃娃2015/10/10Anson.w金刚熊猫娃娃2015/10/10vincentyzw金刚熊猫娃娃2015/10/10路上看到咲金刚熊猫娃娃2015/10/10YumFeiyoung金刚熊猫娃娃2015/10/10狼魂LY辉金刚熊猫娃娃2015/10/10_Dark金刚熊猫娃娃2015/10/10五月雪0金刚熊猫娃娃2015/10/10L等到烟火清凉金刚熊猫娃娃2015/10/10HYB376398金刚熊猫娃娃2015/10/10李大叔驾到金刚熊猫娃娃2015/10/10德国战车金刚熊猫娃娃2015/10/10回家种庄稼金刚熊猫娃娃2015/10/10追杀那只熊:金刚熊猫娃娃2015/10/10zhu*******金刚熊猫娃娃2015/10/10自you自在金刚熊猫娃娃2015/10/10刘海飞金刚熊猫娃娃2015/10/10Aifangert金刚熊猫娃娃2015/10/10秋雨纷飞金刚熊猫娃娃2015/10/10飞_絮金刚熊猫娃娃2015/10/10zwzyc金刚熊猫娃娃2015/10/10林MMM金刚熊猫娃娃2015/10/10Atalei金刚熊猫娃娃2015/10/10wgh222金刚熊猫娃娃2015/10/11荒废了自由金刚熊猫娃娃2015/10/11醉死萌生金刚熊猫娃娃2015/10/11毛亚兴金刚熊猫娃娃2015/10/11bsplin金刚熊猫娃娃2015/10/11xs猴子金刚熊猫娃娃2015/10/11行云之龙金刚熊猫娃娃2015/10/11老煤油关注10年金刚熊猫娃娃2015/10/11夏日魅风金刚熊猫娃娃2015/10/11wii8金刚熊猫娃娃2015/10/11shawlcy金刚熊猫娃娃2015/10/11我不撤退金刚熊猫娃娃2015/10/11Endy_Jay金刚熊猫娃娃2015/10/111天风1金刚熊猫娃娃2015/10/11lingrain金刚熊猫娃娃2015/10/11fay444金刚熊猫娃娃2015/10/11罗成龙07金刚熊猫娃娃2015/10/11无乜缺金刚熊猫娃娃2015/10/11阿木7999金刚熊猫娃娃2015/10/11飞_絮金刚熊猫娃娃2015/10/11Aaron_醒金刚熊猫娃娃2015/10/11陈king金刚熊猫娃娃2015/10/11维震天下金刚熊猫娃娃2015/10/11Agat金刚熊猫娃娃2015/10/11*********金刚熊猫娃娃2015/10/11zbapollo金刚熊猫娃娃2015/10/11O烟雨江南O金刚熊猫娃娃2015/10/11jed_金刚熊猫娃娃2015/10/11rzqlll金刚熊猫娃娃2015/10/11緣來此道非彼道M码2015/10/11CaryWUM码2015/10/11hello_yangM码2015/10/11落血无痕M码2015/10/11戊午天马M码2015/10/11狄威M码2015/10/11高冷萌iM码2015/10/11逆转大势已去M码2015/10/11爽儿...M码2015/10/11十三小师弟M码2015/10/11挚爱binM码2015/10/11骑牛找马M码2015/10/11沧沧1999M码2015/10/11刘小超uM码2015/10/11梦想2020M码2015/10/11尐孑杰M码2015/10/11蘭瑟M码2015/10/11效仿余生丶M码2015/10/11美柚靖M码2015/10/11Xiao喜根M码2015/10/10用户*********M码2015/10/10TheEndsM码2015/10/10redforceM码2015/10/10a*******M码2015/10/10方块森林M码2015/10/10馨馨xM码2015/10/10用户*********M码2015/10/10雨打浮萍泪倾城M码2015/10/10用户********M码2015/10/10ANSYS12M码2015/10/10lilups********M码2015/10/10yyd3250M码2015/10/10小小強M码2015/10/10love*********M码2015/10/10海辛M码2015/10/10七里秋风M码2015/10/9tangyongskyM码2015/10/9路可___M码2015/10/9名字真多好难取M码2015/10/9被啃弯的月亮M码2015/10/9亮剑长空M码2015/10/9♂魅力boyM码2015/10/9古韵筝鸣M码2015/10/9gad_cnM码2015/10/9主上衍安M码2015/10/9Bin氏初级贤M码2015/10/9vaioyfM码2015/10/9zhangguizhuM码2015/10/9转角见到你M码2015/10/9火车怪客eskareM码2015/10/9夜已经深了M码2015/10/9终不济事M码2015/10/9H振祥M码2015/10/8neesonzhaoM码2015/10/8guojie30363M码2015/10/8用户********M码2015/10/8wqvberdaM码2015/10/8用户********M码2015/10/8倾雨漫心M码2015/10/8魑魅魍魉惊本身M码2015/10/8回忆ztM码2015/10/8莳绱丄暧MM码2015/10/8123luohhM码2015/10/8雲先森M码2015/10/8用户********M码2015/10/8花语留芳M码2015/10/8小飞丿o_OM码2015/10/8cladmyM码2015/10/8伯文艺M码2015/10/8沉默的香烟M码2015/10/8枉生jastM码2015/10/8俺是M族M码2015/10/8天地一蜉蝣M码2015/10/8w********M码2015/10/8余轩M码2015/10/8T_mac_糖糖M码2015/10/8贺新M码2015/10/8门生古界M码2015/10/8起风而益M码2015/10/8见朕骑机的时刻M码2015/10/7失乐喵M码2015/10/7sim15M码2015/10/7尐吜渔M码2015/10/7魅911M码2015/10/7TumblingM码2015/10/7喜欢清风M码2015/10/7幻影流风M码2015/10/7凯小龙M码2015/10/7begingoM码2015/10/7徐伤M码2015/10/7qq*******M码2015/10/7佳华流年M码2015/10/7飘洛M码2015/10/7youareaxM码2015/10/7飞翔的寂寞M码2015/10/7梦想伤不起M码2015/10/7puppydoghkM码2015/10/7fastlinM码2015/10/7hhylxcM码2015/10/7haidaofeiM码2015/10/7LesuryeeM码2015/10/7mokaprinceM码2015/10/7zfh3128M码2015/10/6忧郁的蓝色天空M码2015/10/6toatiantM码2015/10/6清水雷明M码2015/10/6落血无痕M码2015/10/6重庆小韩M码2015/10/6jienlM码2015/10/6你是谁0513M码2015/10/6********M码2015/10/6Cyan_DevilM码2015/10/6老虎想猫了M码2015/10/6nevy555M码2015/10/6猴戈M码2015/10/6活着要疯狂M码2015/10/6花自飘零11M码2015/10/6坚持梦想会有奇迹M码2015/10/6Sky苏苏M码2015/10/6quanxiM码2015/10/6kousuidangoM码2015/10/6爱_无言M码2015/10/6FKJJ1985M码2015/10/6小鬼力力.M码2015/10/6羽亦风M码2015/10/6尼克卡卡M码2015/10/5king_88888M码2015/10/5三道杠*好青年M码2015/10/5夢想_LM码2015/10/5未来执法官M码2015/10/5活一天是一天M码2015/10/5初来乍到813M码2015/10/5jonelvM码2015/10/5dragonflyhanM码2015/10/5我是魅蓝M码2015/10/5怎么会呢M码2015/10/5轻轻叩击M码2015/10/5魅呀呀M码2015/10/5择沓M码2015/10/5翔云__追梦M码2015/10/5bqf2M码2015/10/5leishubingM码2015/10/5巨可可M码2015/10/5inourhouseM码2015/10/5hotlogoM码2015/10/5dan********M码2015/10/5|http://bbs.meizu.cn/thread-5750224-1-1.html|2015-10-14
其他媒体|2062445351|difang CN|地方频道 > 滚动读报|ZHO|2015-10-14 14:06:03|上海滩烽烟再起 k3s剑指王座|一次激烈的比赛 一场胜利的狂欢。9月27日 时值万家团圆的中秋佳节 ctcc在上海嘉定烽火重燃。在超级量产组比赛中 东风悦达起亚车队起跑急速突破、转弯行云流水 经过一轮激烈角逐后 小将叶弘历最终力挫群雄 登顶冠军王座。ctcc赛事是梦想的延续 亦是对优秀品质的诠释 东风悦达起亚秉承着“智造经典惠创未来”的经营理念 希望根据中国消费者的喜好持续锻造出更出色的产品 不断给消费者带来更时尚、激情的驾乘体验。|http://difang.gmw.cn/newspaper/2015-10/14/content_109539546.htm|2015-10-14
其他媒体|2064291487|zhidao_baidu|电子数码|ZHO|2015-10-15 13:26:02|东风悦达起亚k3全部费用加一起多少钱|来自：手机知道汽车东风悦达起亚k3全部费用加一起多少钱|http://zhidao.baidu.com/question/874583610649280732.html?fr=qlquick&entry=qb_list_default|2015-10-15
其他媒体|2075149492|zhidao_baidu|全部问题 > 社会民生|ZHO|2015-10-21 17:47:22|东风悦达起亚k3自动挡变速箱r怎么不现视|来自：手机知道汽车东风悦达起亚k3自动挡变速箱r怎么不现视|http://zhidao.baidu.com/question/1606645083602424267.html?fr=qlquick&entry=qb_list_default|2015-10-21
其他媒体|2075167564|zhidao_baidu|东芝|ZHO|2015-10-21 17:58:01|东风悦达起亚k3自动挡变速箱r怎么不现视|来自：手机知道汽车东风悦达起亚k3自动挡变速箱r怎么不现视|http://zhidao.baidu.com/question/1756581186950053508.html?fr=qlquick&entry=qb_list_default|2015-10-21
其他媒体|2075658796|zhidao_baidu|电脑/网络 > 硬件 > 内存|ZHO|2015-10-21 22:53:03|东风悦达起亚k3eco起步好慢|来自：手机知道汽车|http://zhidao.baidu.com/question/1112736334373406259.html?fr=qlquick&entry=qb_list_default|2015-10-21
其他媒体|2178718506|bitauto|易车 > 问答 > 问题分类|ZHO|2015-12-19 20:01:02|起亚k3和本田凌派那个家庭实用些|起亚k3和本田凌派那个家庭实用些     提问者：汽车报价大全**********  分类：  本田  凌派  买车  选车  浏览[6] 来自：汽车报价大全  2015-12-19 18:56  举报   相关车型：凌派 起亚K3|http://ask.bitauto.com/detail/6003299/|2015-12-19
其他媒体|2178950345|difang CN|地方频道 > 滚动读报|ZHO|2015-12-19 23:48:03|2016款吉利新帝豪正式上市|"12月11日 吉利汽车宣布2016款新帝豪正式上市|共推出1.5l和1.3t两种排量9款车型 售价为6.98—10.08万元。2016款吉利新帝豪的推出|不仅体现了帝豪产品品质的不断向上|增配不加价的诚意定价也提高了产品市场竞争力|进一步巩固了帝豪在中国品牌轿车的冠军地位。造型上 2016款吉利新帝豪延续了现款时尚大气、年轻动感的设计风格 并对前脸、车身、尾部等细节处处细节人性化升级。内饰上 新车搭载了全新6向电动调节人机皮质座椅 以酷黑为主色调 全系标配厂家原装脚垫等细节 进一步提升了整车品质。空间上 2016款新帝豪对储物空间进行了多项人性化升级 中控盖板顺应消费者需求改成储物盒设计 中央通道水杯架储物空间拓展等 进一步丰富了车内储物空间。操控方面 2016款吉利新帝豪由英国prodrive（阿斯顿马丁唯一车辆技术合作伙伴）对底盘二次优化 加上美国trw提供的eps电动助力转向 提升了悬挂操纵性与舒适性。动力方面 搭载了吉利自主研发的1.3t和1.5l两款高效绿色节能发动机 匹配六速手动变速器和cvt无级变速器。另外 2016款新帝豪全系车型还能享受3000元节能惠民补贴和购置税减半政策。配置上 全新升级的g-netlink3.0吉利智能车载系统 搭载carplay功能 使用起来更加快捷、方便。安全方面 除1.5mt最低配外 2016款新帝豪全系车型标配新升级的esc车身稳定控制系统 大幅提升安全性能。左小青"|http://difang.gmw.cn/newspaper/2015-12/19/content_110269837.htm|2015-12-19
其他媒体|2180394695|difang CN|地方频道 > 滚动读报|ZHO|2015-12-21 04:20:01|浪漫平安夜与k3暖心出游|圣诞节即将来临 街道上到处呈现出温馨、甜蜜的气息。此时盛装打扮的你 正需要一辆暖心座驾 来感受这个美轮美奂的童话世界。东风悦达起亚k3带着满车的浪漫情怀 伴你感受这欢乐的氛围。k3为你的平安夜打造了暖心的专享空间。k3车身长宽高分别为4600mm、1780mm、1445mm 轴距长达2700mm 带来十分宽敞的内部空间。车舱内 k3运用高档、环保的饰材进行布置 包括具备记忆、加热、通风功能的电动真皮座椅 以及真皮方向盘和门护板、仪表盘等采用的皮包裹设计 让驾乘者感受到了科技魅力所在。另外 凭借n.v.h优化措施 k3还为驾乘者带来了仿佛远离都市般的宁静车舱。（宗合）|http://difang.gmw.cn/newspaper/2015-12/21/content_110284089.htm|2015-12-21
기타|2187705604|315che|行情|ZHO|2015-12-25 13:19:02|起亚K3店内现车充足 购车最高优惠2.2万|　　【上海行情】近日 中国汽车消费网编辑从上海红悦汽车销售服务有限公司了解到 店内起亚K3现车销售 颜色可选 目前购车部分车型可优惠2.20万元。感兴趣的消费者可以进店了解详情 以下是2015款起亚K3的具体的报价表：上海地区起亚4S店最新价格：起亚K3报价表（2015-12-25）车型指导价销售价优惠情况现车情况起亚K3 2015款 1.6L MT GL10.28万8.28万2.0万现车充足起亚K3 2015款 1.6L AT GL11.28万9.28万2.0万现车充足起亚K3 2015款 1.6L AT GLS12.48万10.28万2.2万现车充足起亚K3 2015款 1.6L AT DLX13.18万10.98万2.2万现车充足起亚K3 2015款 1.6L AT Premium14.38万12.18万2.2万现车充足起亚K3 2015款 1.8L AT Premium14.98万12.78万2.2万现车充足中国汽车消费网制表　　起亚K3各地行情信息请关注：http://auto.315che.com/qiyak3/articles__43.htm　　更多同级别车型价格变动信息请关注：http://www.315che.com/hq/　　基本介绍：2015款K3的前中网颜色变更 后保险杠和排气管也经过了重新设计 DLX AT及以上车型配备了椭圆形的镀铬排气管。2015款K3还新增珍珠白这一可选车身颜色。中控面板位置的空调按钮增加镀铬装饰 车内引入了更多软性材料装饰。2015款K3的主要竞争对手还是目前市场上主流的紧凑型轿车 例如现代朗动、本田凌派、雪佛兰科鲁兹等。和竞争对手相比 丰富的配置和个性的造型是吸引不少消费者选择K3的因素。  起亚K3 指导价： 10.28～14.98 万   品牌：起亚图片(共767 张)   配置   车吧   报价   口碑(共133 条)315che.com 　　配置详解：GL配备了主副驾驶座安全气囊、ABS+EBD、多功能方向盘上下调节、行车电脑显示屏、前座中央扶手、前雾灯、大灯高度可调、后视镜电动调节、后视镜加热、手动空调。　　GLS多了日间行车灯、后排杯架、后座中央扶手、座椅高低调节、真皮方向盘、电动天窗、无钥匙启动系统以及选装配置倒车视频影像、真皮座椅、腰部支撑调节、前排座椅电动调节、电动座椅记忆、座椅通风、GPS导航系统、蓝牙/车载电话等。　　DLX在GLS的基础上又多了EBD+EBA+ASR、真皮座椅、后座出风口和温度分区控制。　　Premium作为最高配 新增了后视镜电动折叠、后视镜记忆、氙气大灯、电动座椅记忆、前排座椅加热、座椅通风、前排座椅电动调节、腰部支撑调节、方向盘换挡、定速巡航、胎压监测装置。自动挡还可选装前/后排头部气囊(气帘)。　　注：中国汽车消费网 (www.315che.com) 提供的价格信息为编辑采集的及时信息 价格仅供参考 车市行情天天变 消费者如需购买相关车型 应该尽快与具体经销商电联或当面洽谈。另 文中引用图片和推荐经销商仅为资料信息 与价格信息来源无关。|http://inf.315che.com/n/2015_12/660226/|2015-12-25
其他媒体|2188175549|zhidao_baidu|电脑/网络 > 电脑装机|ZHO|2015-12-25 20:17:02|东风悦达起亚xk3自动档中配大概售价多少钱|汽车东风悦达起亚xk3自动档中配大概售价多少钱|http://zhidao.baidu.com/question/393061427163182725.html?fr=qlquick&entry=qb_list_default|2015-12-25
其他媒体|2216502699|zhidao_baidu|文化/艺术|ZHO|2016-01-11 21:25:01|东风悦达起亚k3油箱多少升|汽车东风悦达起亚k3油箱多少升|http://zhidao.baidu.com/question/1448466591988603380.html?fr=qlquick&entry=qb_list_default|2016-01-11
其他媒体|2244375617|zhidao_baidu|电脑/网络 > 电脑装机|ZHO|2016-01-27 00:16:01|"东风悦达起亚 k3|2015款手动 gl 有日间行车灯吗?"|汽车|http://zhidao.baidu.com/question/265588921927767685.html?fr=qlquick&entry=qb_list_default|2016-01-27
其他媒体|2245493539|youku|时尚|ZHO|2016-01-27 15:11:01|美憬幸感小护士之轮廓注射|小V脸立现的超好评治疗项目！	小V脸立现的超好评治疗项目！隐藏		2小时前 上传|http://v.youku.com/v_show/id_XMTQ1Nzk3NjE0OA==.html|2016-01-27
其他媒体|2246321330|zhidao_baidu|文化/艺术|ZHO|2016-01-27 23:07:31|东风悦达起亚k3买的话还要强制性买平安保险阜阳|阜阳市|http://zhidao.baidu.com/question/1384986375673763620.html?fr=qlquick&entry=qb_list_default|2016-01-27
其他媒体|2252727432|zhidao_baidu|电子数码 > 手机/通讯-手机购买|ZHO|2016-01-31 15:39:02|在长兴买东风悦达起亚k3代款要什么手续|汽车|http://zhidao.baidu.com/question/1670883695748353947.html?fr=qlquick&entry=qb_list_default|2016-01-31
其他媒体|2274534493|zhidao_baidu|电脑/网络|ZHO|2016-02-13 09:42:01|我不知道该选哪款车 以朗动手动领先型对比宝来、k3、英朗、和哈弗h6我该选择哪个 请度友们给点建议|汽车生活以朗动手动领先型对比宝来、和哈弗h6我该选择哪个、k3、英朗 请度友们给点建议我不知道该选哪款车|http://zhidao.baidu.com/question/265788410564983325.html?fr=qlquick&entry=qb_list_default|2016-02-13
기타|2334370189|xcar|导购频道 > 车型海选|ZHO|2016-03-17 05:41:02|销量榜中榜 中国品牌紧凑级轿车争前十|[XCAR 导购 原创]　　前言：近些年 中国品牌汽车的进步是大家有目共睹的 除了中国老牌车企不断壮大外 还有不断涌现的后起之秀。中国品牌在轿车、SUV、MPV等领域多点开花 都取得了骄人的成果。即便SUV现在是热销车型 但三厢轿车在家用车市场依旧有很高的地位。虽说销量并不能完全代表一个产品的好坏 但销量对于消费者来说还是有一定参考价值的。值得一提的是吉利新帝豪在2月份共销售14036辆 成功地挤进轿车销量前十 同时它也是唯一一款进入轿车销量排行榜前十位的中国品牌紧凑级轿车。新帝豪的表现值得称赞 那它的直接竞争对手们表现得又如何？接下来我们将带来三款有能力进入前十的中国品牌紧凑级轿车。    2016年2月轿车销量排名中 中国品牌中仅有吉利新帝豪杀入前十 长安逸动以1049辆的差距紧随其后 虽然上汽荣威360是中国品牌紧凑级销量排名第三位的车型 但销量仅有4483辆 与新帝豪以及逸动的差距较大 但它的实力也绝对不容小觑 假以时日或许也会出现在前十的名单之中。		2016年2月轿车销量排行			排名	车型	2月销量（辆）			1	上汽大众新朗逸	40892			2	一汽-大众速腾	22290			3	上汽通用别克全新英朗	20139			4	上汽大众新桑塔纳	19491			5	一汽丰田卡罗拉	16882			6	一汽-大众捷达	16692			7	长安福特福睿斯	15892			8	上汽通用雪佛兰科鲁兹	15697			9	北京现代朗动	14763			10	吉利帝豪（推荐车型）	14036			12	长安逸动（推荐车型）	12987			20	吉利远景	8379			39	长安悦翔V3	5584			43	吉利金刚	4990			45	长安奔奔	4709			48	上汽荣威360（推荐车型）	4483			49	一汽海马福美来	4361			56	上汽荣威***-****			59	长安悦翔	3530			61	昌河北斗星	3380			爱卡汽车网制表 www.xcar.com.cn	    通过下方推荐车型基本参数表格不难发现 这三款车型的车身尺寸基本处在同一水平。吉利新帝豪车身长度最长 比车身最短的上汽荣威360多出52mm。长安逸动车身高度最高 但也仅比最矮的吉利新帝豪多出31mm。上汽荣威360与长安逸动在车身宽度与轴距方面打成平手 但高度也仅领先新帝豪20mm 轴距也仅多出10mm。		推荐车型基本参数一览表			参数/车型	吉利新帝豪	长安逸动	上汽荣威360			官方指导价格（单位：万元）	6.98-10.08	7.49-11.79	7.59-12.99			长度(单位:mm)	4***-****-****			宽度(单位:mm)	1***-****-****			高度(单位:mm)	1***-****-****			轴距(单位:mm)	2***-****-****			爱卡汽车网制表 www.xcar.com.cn	    推荐车型（一）：吉利新帝豪    售价区间：6.98-10.08万元    车型特点：外形比较时尚且配置相对丰富。    新帝豪造型比较时尚 前进气格栅与两侧自动头灯连为一体 同时头灯内部做了熏黑处理 整体造型比较运动。保险杠两侧嵌入LED日间行车灯 配合内部银色饰条 给人精致的感觉。车身侧面比例比较协调 腰线贯穿车侧 给人修长的感觉。新帝豪的尾部造型比较紧致 细长的镀铬饰条横贯车尾 与尾灯内部灯组相融合。前进气格栅与两侧自动头灯连为一体且头灯内部做了熏黑处理。  新帝豪尾部细长的镀铬饰条横贯车尾并与尾灯内部灯组相融合。    新帝豪的内饰比较简洁 线条也并不复杂。双色四辐方向盘握感比较舒适 同时除时尚型外其余车型方向盘均采用真皮包裹且配备多功能按键。中控台使用撞色设计 下边缘采用色差明显的饰条勾勒 给人年轻时尚的感觉。除时尚型外 其余车型均配备中控彩色大屏 集成G-Netlink3.0车载互联系统。新帝豪的内饰比较简洁 线条也并不复杂。      新帝豪的车身长宽高尺寸为4631mm/1789mm/1470mm 轴距为2650mm。车内的乘坐空间足够日常使用 同时车内的座椅乘坐也比较舒适。新帝豪除时尚型外 其余车型均配备皮革面料座椅 乘坐比较舒适。常规状态下 新帝豪的行李厢容积为680L 同时全系车型后排座椅靠背均支持按比例放倒。车内的储物空间比较丰富 实用性较高。车内的乘坐空间足够日常使用 同时车内的座椅乘坐也比较舒适。      吉利新帝豪拥有1.3T和1.5L两款发动机 1.3T发动机最大功率为98kW（133Ps）/5500rpm 峰值扭矩为185Nm/****-****rpm 传动系统匹配6挡手动或CVT无级变速箱 工信部公布的手动挡车型综合油耗为5.7L/100km 自动挡车型综合油耗为5.9L/100km。1.5L发动机最大功率为80kW（109Ps）/6000rpm 峰值扭矩为140Nm/4400rpm 传动系统匹配5挡手动或CVT无级变速箱 工信部公布的手动挡车型综合油耗为5.7L/100km 自动挡车型综合油耗为5.9L/100km。悬挂方面 新帝豪采用前麦弗逊式独立悬挂后扭力梁式非独立悬挂的组合。吉利新帝豪拥有1.3T和1.5L两款发动机。1.3T匹配6挡手动或CVT变速箱 1.5L匹配5挡手动或CVT变速箱。新帝豪采用前麦弗逊式独立悬挂后扭力梁式非独立悬挂的组合。    通过2月份销量统计表我们发现 吉利有多款车型都取得了不错的销量 这也间接证明了吉利是在用心造车 吉利汽车也被越来越多的消费者接受 作为目前唯一一款销量挤进前十的中国品牌轿车 新帝豪的实力还是值得肯定的。|http://newcar.xcar.com.cn/201603/news_1917436_1.html|2016-03-17
其他媒体|2334407678|youku|生活|ZHO|2016-03-17 06:40:02|监控实拍：起亚无视大货车 高速野蛮超车 比...|视频: 监控实拍：起亚无视大货车 高速野蛮超车 比亚迪唐吓尿了...|http://v.youku.com/v_show/id_XMTUwMTk3MDYzMg==.html|2016-03-17
其他媒体|2334513728|bitauto|易车 > 问答 > 问题分类|ZHO|2016-03-17 08:43:01|"卡罗拉 朗逸 k3|英朗 宝来 h2 雷凌 朗动 新克鲁兹轩"|"卡罗拉 朗逸 k3|英朗 宝来 h2 雷凌 朗动 新克鲁兹轩     提问者：YCAPP160311C6U9E  分类：  起亚  K3  其他  浏览[12] 来自：易车手机客户端  2016-03-17 07:21  举报   卡罗拉 朗逸 k3|英朗 宝来 h2 雷凌 朗动 新克鲁兹轩逸。哪个好 给个理由和配置 裸车不超12万谢谢了。我好迷茫"|http://ask.bitauto.com/detail/6311923/|2016-03-17
其他媒体|2334513732|bitauto|易车 > 问答 > 问题分类|ZHO|2016-03-17 08:43:01|"#帮我选车# 卡罗拉 朗逸 k3|英朗 宝来 h2 雷凌 朗"|"#帮我选车# 卡罗拉 朗逸 k3|英朗 宝来 h2 雷凌 朗     提问者：YCAPP160311C6U9E  分类：  起亚  K3  买车  选车  浏览[8] 来自：易车手机客户端  2016-03-17 07:21  举报   #帮我选车# 卡罗拉 朗逸 k3|英朗 宝来 h2 雷凌 朗动 新克鲁兹轩逸。哪个好 给个理由和配置 裸车不超12万谢谢了。我好迷茫"|http://ask.bitauto.com/detail/6311925/|2016-03-17
各大媒体|2334887250|qc188|主题导购 > 多功能/其他|ZHO|2016-03-17 12:42:01|有能力进入前十 三款中国品牌紧凑车型|　　前言：近些年 中国品牌汽车的进步是大家有目共睹的 除了中国老牌车企不断壮大外 还有不断涌现的后起之秀。中国品牌在轿车、suv、MPV等领域多点开花 都取得了骄人的成果。即便SUV现在是热销车型 但三厢轿车在家用车市场依旧有很高的地位。虽说销量并不能完全代表一个产品的好坏 但销量对于消费者来说还是有一定参考价值的。值得一提的是吉利新帝豪在2月份共销售14036辆 成功地挤进轿车销量前十 同时它也是唯一一款进入轿车销量排行榜前十位的中国品牌紧凑级轿车。新帝豪的表现值得称赞 那它的直接竞争对手们表现得又如何？接下来我们将带来三款有能力进入前十的中国品牌紧凑级轿车。    2016年2月轿车销量排名中 中国品牌中仅有吉利新帝豪杀入前十 长安逸动以1049辆的差距紧随其后 虽然上汽荣威360是中国品牌紧凑级销量排名第三位的车型 但销量仅有4483辆 与新帝豪以及逸动的差距较大 但它的实力也绝对不容小觑 假以时日或许也会出现在前十的名单之中。2016年2月轿车销量排行排名车型2月销量（辆）1上汽大众新朗逸408922一汽-大众速腾222903上汽通用别克全新英朗201394上汽大众新桑塔纳194915一汽丰田卡罗拉168826一汽-大众捷达166927长安福特福睿斯158928上汽通用雪佛兰科鲁兹156979北京现代朗动1476310吉利帝豪（推荐车型）1403612长安逸动（推荐车型）1298720吉利远景837939长安悦翔V3558443吉利金刚499045长安奔奔470948上汽荣威360（推荐车型）448349一汽海马福美来436156上汽荣威***-****59长安悦翔353061昌河北斗星3380    通过下方推荐车型基本参数表格不难发现 这三款车型的车身尺寸基本处在同一水平。吉利新帝豪车身长度最长 比车身最短的上汽荣威360多出52mm。长安逸动车身高度最高 但也仅比最矮的吉利新帝豪多出31mm。上汽荣威360与长安逸动在车身宽度与轴距方面打成平手 但高度也仅领先新帝豪20mm 轴距也仅多出10mm。推荐车型基本参数一览表参数/车型吉利新帝豪长安逸动上汽荣威360官方指导价格（单位：万元）6.98-10.087.49-11.797.59-12.99长度(单位:mm)4***-****-****宽度(单位:mm)1***-****-****高度(单位:mm)1***-****-****轴距(单位:mm)2***-****-****    推荐车型（一）：吉利新帝豪    售价区间：6.98-10.08万元    车型特点：外形比较时尚且配置相对丰富。    新帝豪造型比较时尚 前进气格栅与两侧自动头灯连为一体 同时头灯内部做了熏黑处理 整体造型比较运动。保险杠两侧嵌入LED日间行车灯 配合内部银色饰条 给人精致的感觉。车身侧面比例比较协调 腰线贯穿车侧 给人修长的感觉。新帝豪的尾部造型比较紧致 细长的镀铬饰条横贯车尾 与尾灯内部灯组相融合。前进气格栅与两侧自动头灯连为一体且头灯内部做了熏黑处理。  新帝豪尾部细长的镀铬饰条横贯车尾并与尾灯内部灯组相融合。    新帝豪的内饰比较简洁 线条也并不复杂。双色四辐方向盘握感比较舒适 同时除时尚型外其余车型方向盘均采用真皮包裹且配备多功能按键。中控台使用撞色设计 下边缘采用色差明显的饰条勾勒 给人年轻时尚的感觉。除时尚型外 其余车型均配备中控彩色大屏 集成G-Netlink3.0车载互联系统。新帝豪的内饰比较简洁 线条也并不复杂。      新帝豪的车身长宽高尺寸为4631mm/1789mm/1470mm 轴距为2650mm。车内的乘坐空间足够日常使用 同时车内的座椅乘坐也比较舒适。新帝豪除时尚型外 其余车型均配备皮革面料座椅 乘坐比较舒适。常规状态下 新帝豪的行李厢容积为680L 同时全系车型后排座椅靠背均支持按比例放倒。车内的储物空间比较丰富 实用性较高。车内的乘坐空间足够日常使用 同时车内的座椅乘坐也比较舒适。      吉利新帝豪拥有1.3T和1.5L两款发动机 1.3T发动机最大功率为98kW（133Ps）/5500rpm 峰值扭矩为185Nm/****-****rpm 传动系统匹配6挡手动或CVT无级变速箱 工信部公布的手动挡车型综合油耗为5.7L/100km 自动挡车型综合油耗为5.9L/100km。1.5L发动机最大功率为80kW（109Ps）/6000rpm 峰值扭矩为140Nm/4400rpm 传动系统匹配5挡手动或CVT无级变速箱 工信部公布的手动挡车型综合油耗为5.7L/100km 自动挡车型综合油耗为5.9L/100km。悬挂方面 新帝豪采用前麦弗逊式独立悬挂后扭力梁式非独立悬挂的组合。吉利新帝豪拥有1.3T和1.5L两款发动机。1.3T匹配6挡手动或CVT变速箱 1.5L匹配5挡手动或CVT变速箱。新帝豪采用前麦弗逊式独立悬挂后扭力梁式非独立悬挂的组合。    通过2月份销量统计表我们发现 吉利有多款车型都取得了不错的销量 这也间接证明了吉利是在用心造车 吉利汽车也被越来越多的消费者接受 作为目前唯一一款销量挤进前十的中国品牌轿车 新帝豪的实力还是值得肯定的。  [1] [2] [3] [下一页] 大家都在关注这些导购：6万左右两厢车 4万左右的三厢车 6万元家用车 12万以内的车 10万元合资suv 100万左右的车 10万以下两厢车|http://www.qc188.com/ztdg/201603/20745.html|2016-03-17
其他媒体|2336033104|bitauto|汽车行情 RSS|ZHO|2016-03-18 00:24:02|【长安CS75深圳官方车友会】DSA深圳车友会版及最新地图资|"生 命 不 息   折 腾 不 止 ！ ！ ！在国内的CS75车友中 绝对多数的人对CS75的做工 用料及设计等各方面 都是一致的好评 但是导航却又是大家一致的吐槽点 当然 这导航也不是一无是处 大神级的专业电子高手攀枝花【神秘人】的观点 用料 做工和配置都很棒 大家都想不明白为啥只用4G的内存芯片 再整个阉割了大量详地图数据的地图 变成了神一般的导航 可以不停的让你转圈圈 可以让你上天入地无所不能 可以让车开到海里去 还能开出来。世上无难事 只怕有心人 经常全国各地一帮子爱折腾的家伙夜以继日的鼓捣 发挥大家各自的长处 相互交流学习 溶合等等 总之花费了大家大量的心血 并经常大量的改装之后 总结经验慢慢的形成了大体固定的改装方案。硬件方面 在最早的南京金陵极速车友会 【老虾】 大神的芯片脚焊线外置TF卡后 大体形成如下两个被广泛采用改装方案：1.攀枝花神秘人针对有电子基础车友的方案 杜邦线+卡槽 直接在主板上预留的卡槽位上焊线 第四脚跳线到元件C220处 卡槽放在导航右侧空出来的按键处。特点 稳定 读不到卡的机率极低 但是按键开孔是个技术活 建议车友们直接把卡槽粘机器外 简单省事。2.深圳车友会小廖原创针对菜鸟车友的的方案 主板焊翻盖式卡槽+20CM延长线 压敏电阻FB2移到FB10处 卡槽粘机器外的方案 所有部件均可网上采购 然后找修手机的师傅 按图操作 自己拷贝软件就OK了。特点 配件易采购 自己少动手 但是读不到卡 黑屏白线的机率略高 黑屏白线的原因就是没读到TF卡 大家检查一下 找到原因就行了。 我们的车标易车大旗 现在小廖的TF卡槽基本是这样放的 线短稳定 藏起来更美观 一年更新一次 拆下猪耳朵就行了。在此增加一个困扰很多人的问题的改解方案：黄星不定位的问题。黄星不定位 说明机器搜星和硬件都是正常的 问题产生的原因是干扰 车内外来的干扰设备极少 经过数次查找 最后发现是射频发生器产生的干扰。射频发生器的位置在主驾遮阳板后 拆下顶灯 左边的插头插着的就是那个东东。解决方案如下：部份车辆是外置后装机第一次导航不定位 请点开导航软件中的GPS卫星状态 如果出现黄星 启动发动机后拆下顶灯 拔掉射频发生器插头 让导航定位后再插上 如果马上掉星 请辅以收音机搜台模式 搜台一次 并重新启动 如果正常搜星定位 则问题解决；如果重复数次依黄星不定位 则需要去4S保修更换射频发生器了。注：拔下射频发生器以后 车辆是无法接收遥控钥匙的信号 不解码发动机的电子防盗系统是无法启动发机的 烦请注意！！下面的话可能会招来鄙视和骂声一遍：你个死胖纸 不吹水你会死啊！！！但我还是要说 黄星不定位是射频发生器的干扰 CS75深圳小廖是国内CS75导航改装圈中第一个找到根本原因所在的死胖纸！！ 黄星不定位是这个样子的。软件方面在经过最早的DSA+地图 再到【萌萌哒抠脚大汉】的一机多图 一机多图简化版 再到车友【Lee】针对网络软件改进的一机多图WIN8版等等。大家为了CS75导航 也因为各自的爱好 花费大量心血 做了大量的贡献 不断的给全国的CS75车友以惊喜 我们应当感谢他们 此处因有鲜花和掌声。当然 我们的折腾行为 在16年会慢慢的部分划上句号 除了之前车主需要继续折腾外 从16款CS75开始 车载导航换成了内存16G的安卓机 经过小廖实车测试 16款导航的屏幕更加细腻 显示分辨率有所提升 反应速度敏捷 地图数据也很详细 最大的改善来自于导航路径的选择更为人性化。只是对于大部分用习惯了凯立德导航的车友们 需要一个智暂的适应过程。--------------------------------------------------------------------------------------------------------------------------------------------------------------------- 硬件差不多了 软件因为不是专用程序 车友们都是要边测试变修改 使用中发现问题目后再修改甚至推倒重来 不断的改进优化 争取让软件和我们的导航更匹配 运行更稳定 更漂亮 以及需要不断更新的地图资源。最近很长一段时间 副会长老廖同志都是悄无声息 问他原因 他才透露 一直在黙默的改写和测试导航主界面软件及地图资源。忙碌中接到他的电话 软件测试完全 可以装车并发布了 带着激动的心情 开着我的骚红小7出发了！！干嘛呢？？？当然是去拿软件。 对你爱 爱 爱不完副会长   002福永-老廖    感谢老廖 一直以来在背后黙黙的支持和付出！ 今天给大家带来的是【长安CS75深圳车友会】002副会长老廖经过一两个月 利用工作之余的时间 花费大量精力改写的程序【善领DSA P57深圳车友会2.5版】、【善领DSA深圳车友会卡拉OK版】、【善领DSA P56深圳车友会1.0版】【一机多图深圳车友会5.2专版】 【一机多图WIN8版】以及经过无数次实测 针对75导航做了适应性数据修改 以及使用中的操作注意事项 2016年3月最新的地图资源。 本帖所有资料源仅作为交流使用 作死有风险 动手需谨慎 由些带来的后果 请自负。以下为相关资源及说明图片： 【善领DSA P57深圳车友会2.5版】https://yunpan.cn/cY6v7vEMSvDpX  访问密码 bab9   晚上的界面  【善领DSA深圳车友会卡拉OK版】https://yunpan.cn/cYMUIXtTEzevd  访问密码 15ca 善领DSA P56深圳车友会1.0版】https://yunpan.cn/cY62sjtI49GRA  访问密码 315d    1.0版 晚上的界面 来自车友【Lee】的 【一机多图WIN8版】版本https://yunpan.cn/cYERk387LFwJv  访问密码 fc18  一机多图WIN8版简化界面  【一机多图深圳车友会5.2专版】https://yunpan.cn/cYMzg6axyyxcs  访问密码 b927 老廖同志根据网络原程序修改的【WIN8一机多图深圳车友会5.1版】https://yunpan.cn/cYY26zcPr5s3Y  访问密码 7920我们将对稳定性和功能做进一步的优化和简化以下为地图资源本资源所有地图资源均来自于网络论坛：我爱GPS GPS之窗 感谢各位大神的力作 本资源只能作为车友之间的交流使用 不得作为商业用途 特此说明。本资源所有地图软件 均经过【长安CS75深圳官方车友会】副会长老廖同志的实测 暂未发现问题 如有问题 烦请和【长安CS75深圳官方车友会】（QQ群号：425338O41）联系 谢谢！！A 地图版本号凯立德（自适应版）：凯立德冬季正式版主程序C3261-C7M10-3821J0Q凯立德（端口版）：凯立德冬季正式版主程序C3261-C7M10-3821J0Q图吧： 83139+NBF12美行： ***.***.***.***CA（Z17）道道通：版本本号:RT-H1A-22AW-K高德： V31（主要用于同步导航系统时间）地图文件中的 凯立德3821（自适应版）、图吧、美行、道道通 均为自适应端口 无需改数据。直接解压后请将文件夹放在TF卡里 并一机多图 DSA和其他地图文件并列 详情见安装目录参考样图。凯立德3821（端口版）和高德V31|在DSA+地图包的模式引领下 端口为：COM8 比特率：9600 ；在一机多图引领下|端口为：COM1 比物率：9600注意：高德在一机多图下 只能选在界面直接进入和DSA引领下进入二选一 不支持都可以进入。界面直接进入 请用端口工具将端口修改为：COM1比特率：9600 DSA进入端口：COM8 比特率：9600凯立德3821（自适应版） 同样为一机多图和DSA引领二先一。在第一次导航进入地图时 会自动适配车机数据 并产生配置文件保存 所以 第一次开机时在一机多图下直接进入的 以后都只能在一机多图下进入 DSA下无法定位；第一次在DSA导航路径下进入的 以后都只能从DSA导航路径下进入。装有凯立德3821（自适应版）的TF卡 只能在第一次试机的导航上用 换到其他导航时 需要重新拷贝地图文件。凯立德3821（端口版）则与之前的操作方式一样 可以实现一机多图下 界面和DSA均可进入 请用端口工具将端口修改为：COM1比特率：9600 DSA进入端口：COM8 比特率：9600 一机多图下DSA的凯立德导航引导路径：App/XSS/KLD.EXE凯立德c3261-c7m10-3821（sp1）下载主程序加入地图包文件构成凯立德大小6.72 G 这不是3D版 因为是自适配端口 所以上机后先不能运行 如果在DSA里运行请先设置好路径等待DSA搜星正常后再点击凯立德 适配完成后就能在DSA正常运行 如果在一机多图里运行（想独立运行）操作方法和上面一样 适配成功后一机多图界面就可以运行（只能二选一 要么DSA里运行 要么一机多图界面运行）。注：经测试 凯立德3821（自适应版）运行速度度更快；凯立德3821（3D端口版）运行速度相对较慢一些。 一机多图TF卡目录下文件夹的参考图   DSA+多地图TF卡目录下文件夹的参考图   凯立德（自适应版）：凯立德冬季正式版主程序C3261-C7M10-3821J0Q https://yunpan.cn/cYMpshfCnwBap  访问密码 3375凯立德（3D端口版）：凯立德冬季正式版主程序C3261-C7M10-3821J0Qhttps://yunpan.cn/cYMpKuSpgek4J  访问密码 b943凯立德（3D端口版）端口修改工具https://yunpan.cn/cYMpVcVdkzgTg  访问密码 ca30 图吧：  83139+NBF12https://yunpan.cn/cYMpLHDrZqTYP  访问密码 d32d 美行：  ***.***.***.***CA（Z17）https://yunpan.cn/cYMpuyKIKdpN8  访问密码 4a44道道通：版本本号:RT-H1A-22AW-Khttps://yunpan.cn/cYMpxL7mszd48  访问密码 d80d 高德： V31（主要用于同步导航系统时间）https://yunpan.cn/cYMpq57QUBbQp 访问密码 9b2a高德端口修改工具：https://yunpan.cn/cYMpW83GhAXXB 访问密码 c786WIN CE5.0游戏包：https://yunpan.cn/cYMppMtHAWFny 访问密码 990eWIN CE5.0游戏包 通过DSA引领时 需要通过导航路径设定指引运行 才可以使用。在一机多图中使用时 放到TF卡目录下 点击界面上的游戏进入使用。导航各种路径引导的配置文件（因需选用 仅供参考：https://yunpan.cn/cY6vaF7RdUImL 访问密码 a52c  再 次 声 明：本帖所有资料源仅作为交流使用 作死有风险 动手需谨慎 由些带来的后果 请自负。本资源所有地图资源均来自于网络论坛：我爱GPS GPS之窗 感谢各位大神的力作 本资源只能作为车友之间的交流使用 不得作为商业用途 特此说明。愿大家：人 长 久  车 长 安 ！！深圳周边 喜欢和想了解CS75的朋友 欢迎加入我们的预备群：【深圳CS75官方车友会预备群】（QQ群号：*********） 我们将用大家真实的使用体验与心得 为你解答与CS75相关的问题！！【长安CS75深圳官方车友会】（QQ群号：*********） 深圳地区【唯一】【长安汽车】【厂家认证】的CS75官方车友会！深圳福利最好、最给力的纯75车主的车友会 期待CS75车主您的加入 我们将用富有自己特色的生活方式 丰富的改装经验及资源、丰厚的售后福利及大量的自驾游和交流活动 在和75相伴的日子里 活出不一样的精彩！     0"|http://bitauto.feedsportal.com/c/33450/f/584188/s/4e555d39/sc/33/l/0Lbaa0Bbitauto0N0Cchangancs750Cthread0E88163290Bhtml/story01.htm|2016-03-18
기타|2336657217|163_bbs|网易新闻论坛-社会万象|ZHO|2016-03-18 11:00:01|被杨幂一手带大的迪丽热巴真的要把杨幂...|一手带大的迪丽热巴 颜值要开始追赶了  无论哪个角度都美啊  可爱的胖迪  “痴呆”少女既视感啊  美如画的侧面  身材很棒啊！~  真的是要替代杨幂成为最新小花啊！~ http://www.aspcms.com/cdjk/hys69/***************74.html http://whjk.zznews.cn/gytu/***************29.html http://top.123cha.com/fr95q/***************81.html http://www.47.etobq.top/ http://top.123cha.com/fghgf8tr/***************00.html http://yunjk.123cha.com/bfbf14/***************01.html http://top.123cha.com/cvhdre3/***************50.html http://www.aspcms.com/cdjk/wwqrt/***************73.html http://2013diebian.*******.com/d14/***************68.html http://whjk.zznews.cn/swer/***************15.html http://j3x.w34o.hkfrx.top/ http://www.rpc.urbxn.cn/ http://yunjk.123cha.com/cghy/***************89.html http://www.aspcms.com/cdjk/wwqrt/***************43.html http://kxw.o2fi.mrufm.top/ http://ep5.ccwujing.website/ http://top.123cha.com/cvhdre3/***************88.html http://ycjk.ltaaa.com/y0u/***************32.html http://kc62.x6cg.sxcxtz.cricket/ http://top.123cha.com/y2d9s/***************78.html http://ycjk.ltaaa.com/y0u/***************01.html http://top.123cha.com/fr95q/***************99.html http://whjk.zznews.cn/fgfhf18/***************59.html http://whjk.zznews.cn/gytu/***************56.html http://www.o2hw.byxyf.xyz/ http://yunjk.123cha.com/fgfbfb65/***************54.html http://2013diebian.*******.com/c14/***************19.html http://ehg.m137.52fkw.cn/ http://3im.lxo5.shenbingke120.cn/ http://ycjk.ltaaa.com/lin0/***************22.html http://www.3wbu.mapgd.date/ http://www.aspcms.com/cdjk/vbhm/***************10.html http://whjk.zznews.cn/dvfbg15/***************46.html http://yunjk.123cha.com/cghy/***************91.html http://whjk.zznews.cn/fgfhf18/***************96.html http://www.aspcms.com/cdjk/gt0sw/***************90.html http://www.s7c.vjehn.cn/ http://yunjk.123cha.com/fr36q/***************31.html http://www.aspcms.com/cdjk/dvfdvbf45/***************86.html http://top.123cha.com/y2d9s/***************23.html http://njd.mrg8.btexr.cn/ http://vb2.e1x6.flxfd04.cn/ http://bmld.ack1.bzhvcj4.cn/ http://qvt.xtqo.tnaz800.cn/ http://top.123cha.com/cvhdre3/***************54.html http://top.123cha.com/fghgf8tr/***************33.html http://www.aspcms.com/cdjk/vbhm/***************99.html http://whjk.zznews.cn/fgfhf18/***************74.html http://2013diebian.*******.com/g15/***************88.html http://www.aspcms.com/cdjk/vbhm/***************67.html http://www.aspcms.com/cdjk/dvfdvbf45/***************63.html http://top.123cha.com/cvhdre3/***************06.html http://www.aspcms.com/cdjk/wwqrt/***************14.html http://whjk.zznews.cn/gytu/***************76.html http://whjk.zznews.cn/ups0w/***************28.html http://ycjk.ltaaa.com/r10/***************84.html http://5z3.24us.eaear.top/ http://top.123cha.com/fghgf8tr/***************24.html http://www.aspcms.com/cdjk/hys69/***************21.html http://www.aspcms.com/cdjk/dvfdvbf45/***************29.html http://yunjk.123cha.com/fgfbfb65/***************05.html http://mafj.uyg7.eigrzm.date/ http://n3m.x4jr.pwtkcj1.cn/ http://www.9kq.afygi.cn/ http://xnqj.nd4.xhavs.xyz/ http://top.123cha.com/vy30e/***************04.html http://madr.n57.pgkdz.date/ http://www.aspcms.com/cdjk/gtq6s/***************97.html http://top.123cha.com/fr95q/***************83.html http://0yr.3rmn.521jk.cn/ http://whjk.zznews.cn/gytu/***************01.html http://2013diebian.*******.com/mv4/***************24.html http://2013diebian.*******.com/d14/***************53.html http://www.aspcms.com/cdjk/wwqrt/***************82.html http://www.7dlj.nuxye.xyz/ http://nf4w.0ek.ruknu.top/ http://www.aspcms.com/cdjk/hys69/***************53.html http://whjk.zznews.cn/swer/***************08.html http://y9ef.0pf.btexr.cn/ http://whjk.zznews.cn/gytu/***************81.html http://yunjk.123cha.com/fgfbfb65/***************88.html http://2013diebian.*******.com/c14/***************13.html http://top.123cha.com/fghgf8tr/***************90.html http://i5k.n823.udltv.cn/ http://www.aspcms.com/cdjk/wwqrt/***************16.html http://ycjk.ltaaa.com/y0u/***************60.html http://whjk.zznews.cn/gytu/***************75.html http://7i5.xe3y.wulis.cn/ http://a05o.vw6.avavm.top/ http://r0qm.dvo4.ccfk120.cn/ http://2013diebian.*******.com/c60/***************29.html http://2013diebian.*******.com/g15/***************45.html http://www.tf.texwyf.cricket/ http://whjk.zznews.cn/swer/***************08.html http://ycjk.ltaaa.com/r10/***************69.html http://yunjk.123cha.com/bfbf14/***************84.html http://www.rwv.bwjsb.xyz/ http://www.8cdu.sbkrg.xyz/ http://www.y7xb.wuhanht.date/ http://Yv.ccygyy.cn/ http://2013diebian.*******.com/c60/***************46.html http://ekq7.lcy.afygi.cn/ http://2013diebian.*******.com/c60/***************67.html http://ycjk.ltaaa.com/e79/***************74.html http://yunjk.123cha.com/hygf/***************39.html http://2013diebian.*******.com/c60/***************61.html http://ido0.vdkt.dbqtve.cricket/ http://ycjk.ltaaa.com/y0u/***************23.html http://yunjk.123cha.com/hygf/***************43.html http://whjk.zznews.cn/hy29a/***************85.html http://8a1.2yc3.shengbingke120.cn/ http://top.123cha.com/fghgf8tr/***************58.html http://yunjk.123cha.com/cghy/***************89.html http://w9n.gf0a.********.cn/ http://yunjk.123cha.com/fgfbfb65/***************93.html http://2013diebian.*******.com/c14/***************53.html http://whjk.zznews.cn/gytu/***************15.html http://xmof05.sbk39.website/ http://6g49.yump.wjsk1199.website/ http://vehd.x1j.wkweo.cc/ http://yunjk.123cha.com/fgfbfb65/***************86.html http://yunjk.123cha.com/hygf/***************44.html http://0v4w.4xnp.rlgwvx.cricket/ http://mgd.shenbing120.cn/ http://zhoj.nhx.pbcza.cn/ http://top.123cha.com/y2d9s/***************59.html http://www.sa0c.bwjsb.xyz/ http://www.q51.qumxz.date/ http://ycjk.ltaaa.com/r10/***************55.html http://whjk.zznews.cn/hy29a/***************29.html http://sxz.7o25.0431wjyy.cn/ http://top.123cha.com/cvhdre3/***************17.html http://www.aspcms.com/cdjk/gtq6s/***************49.html http://www.7re.unbmq.xyz/ http://2013diebian.*******.com/c14/***************51.html http://whjk.zznews.cn/gytu/***************03.html http://ycjk.ltaaa.com/r10/***************87.html http://whjk.zznews.cn/gytu/***************63.html http://2013diebian.*******.com/d14/***************42.html http://ycjk.ltaaa.com/c10/***************23.html http://keh.1uxc.********.cn/ http://top.123cha.com/fr95q/***************72.html http://ozpa.ud5.sbkrg.xyz/ http://www.empd.hkfrx.top/ http://whjk.zznews.cn/fgfhf18/***************12.html http://egz.shenneike120.cn/ http://whjk.zznews.cn/fgfhf18/***************57.html http://www.yx30.afygi.cn/ http://2013diebian.*******.com/g4i/***************14.html http://ycjk.ltaaa.com/e79/***************34.html http://lqif.vxoc.208fukew.cn/ http://qbv.bjfu.johzsy.cricket/ http://www.aspcms.com/cdjk/gt0sw/***************72.html http://w3h.ipjxzq.cricket/ http://www.s83.bivfy.date/ http://www.yif.tmjzk.xyz/ http://whjk.zznews.cn/gytu/***************91.html http://top.123cha.com/vy30e/***************73.html http://ejr.24ik.dbbyby.cn/ http://1od2.i7r1.120girl.cn/ http://2013diebian.*******.com/c14/***************98.html http://08v.wulis.cn/ http://www.aspcms.com/cdjk/gt0sw/***************93.html http://www.aspcms.com/cdjk/gt0sw/***************54.html http://whjk.zznews.cn/swer/***************13.html http://www.aspcms.com/cdjk/dvfdvbf45/***************87.html http://1ebu.9me.eaear.top/ http://top.123cha.com/cvhdre3/***************52.html http://2013diebian.*******.com/c60/***************43.html http://h0w6.n7jb.wulis.cn/ http://qi6.ce0y.wvexk.top/ http://fqyg10.skdmc.cn/ http://whjk.zznews.cn/gytu/***************70.html http://9kx.qmdc.cchmfk.cn/ http://2013diebian.*******.com/mv4/***************52.html http://top.123cha.com/cvhdre3/***************04.html http://yunjk.123cha.com/cghy/***************58.html http://q0h.jv9x.cznsu.cn/ http://www.aspcms.com/cdjk/hys69/***************48.html http://********.shenbing120.website/ http://www.2na.gbdcy.xyz/ http://k5l.b0v1.pbcza.cn/ http://octu.9vmu.ccyc120.cn/ http://vmy.3qkm.ccfuke120.cn/|http://bbs.news.163.com/bbs/society/602605562.html|2016-03-18
其他媒体|2336679087|zhidao_baidu|生活 > 购物|ZHO|2016-03-18 11:14:01|东风悦达起亚k3经济行大概多少钱|汽车东风悦达起亚k3经济行大概多少钱|http://zhidao.baidu.com/question/2077162483582107588.html?fr=qlquick&entry=qb_list_default|2016-03-18
其他媒体|2337718483|bitauto|易车 > 问答 > 问题分类|ZHO|2016-03-18 22:14:03|哈佛h2 现代朗动 起亚k3 手动中配的|哈佛h2 现代朗动 起亚k3 手动中配的     提问者：汽车报价大全********  分类：  哈弗  哈弗H2  买车  选车  浏览[6] 来自：汽车报价大全  2016-03-18 21:08  举报   相关车型：哈弗H2 朗动 起亚K3|http://ask.bitauto.com/detail/6318993/|2016-03-18
기타|2376316888|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:02:02|爪 狠狠向其中一只蛇女抓去 |弗兰德惊慌失措的跌下山坡 没等他立足 便死命召唤变异兽向他靠拢 此时众人已到他头顶之上 继续几十枚黏胶炮弹向他们射过来 这次蛇女没敢让那东西粘上自己的护罩 喷出轻易不肯动用的冰蓝寒气将其冻成冰球 接着又有兽化战士背着超新星做人肉炸弹疯狂向下冲来 吓得弗兰德屁滚尿流 恨不能分裂思维 再找一个分身躲过这一劫难 好在他身边的蛇女拥有大型圣魂器 乍然释放出数百米毁灭红光 将飞过来的兽化战士尽皆毁灭。            若不是弗兰德一开始就被吓破了胆子 蛇女们也不是没有一战之力 弗兰德一门心思想要冲进大盐湖 圣魂器的红光乍现既逝 一直被厄俄斯保护好好的迪莉娅主动冲出来 兽化战士只剩下不到二十个 他们不准备白白消耗这些炮灰 面对蛇女的圣魂器 大多数进化者都无能为力 从没有在其他人面前出过手的迪莉娅 一出手就让其他人惊惧不已。            就见迪莉娅小手一挥 一道细长的阴影从她的身上扩展出来快速放大 初时阴影只有五道细细小条 瞬间扩大无数倍 犹如百米龙http://www.pe6.0431rl.cn/    http://www.xsu.0431wjyy.cn/    http://www.hwk.120girl.cn/    http://www.78u.120shenbingke.cn/    http://www.y6t.120shenneike.cn/    http://www.gmt.120szbyy.cn/    http://www.gdf.120wjyy39.cn/    http://www.uaw.208fukew.cn/    http://www.3dg.521jk.cn/    http://www.3i7.52fkw.cn/    http://www.96f.********.cn/    http://www.54y.********.cn/    http://www.g39.********.cn/    http://www.1uc.********.cn/    http://www.0b3.********.cn/    http://www.xqp.********.cn/    http://www.t47.********.cn/    http://www.k0t.********.cn/    http://www.b62.asqnf.cn/    http://www.r89.buyun365.cn/    http://www.q8k.bzhvcj4.cn/    http://www.b78.cc516.cn/    http://www.et5.ccby120.cn/    http://www.9kq.ccbyby.cn/    http://www.ojw.ccfk120.cn/    http://www.w76.ccfkyy.cn/    http://www.m6w.ccfkyy120.cn/    http://www.ftk.ccfuke.cn/    http://www.w53.ccfuke120.cn/    http://www.qn8.cchmfk.cn/    http://www.ceo.ccmly120.cn/    http://www.jrw.ccrenliu.cn/    http://www.7ek.ccrl120.cn/    http://www.4wp.ccrlyy.cn/    http://www.yde.ccrsfk.cn/    http://www.lnu.ccsfuchan.cn/    http://www.sod.ccshenbing120.cn/    http://www.yz9.ccshenbing39.cn/    http://www.toq.ccszbyy120.cn/    http://www.9vp.ccwtrl.cn/    http://www.ozy.ccxhfk.cn/    http://www.8m6.ccyc120.cn/    http://www.qyg.ccyg120.cn/    http://www.3oh.ccygfk.cn/    http://www.i21.ccygfk120.cn/    http://www.va4.ccygyy.cn/    http://www.xq8.ccygyy120.cn/    http://www.ncy.dbbyby.cn/    http://www.6pg.dslr120.cn/    http://www.6fm.eapaz36.cn/    http://www.t2k.fkylw.cn/    http://www.5pc.fkzx120.cn/    http://www.j86.flxfd04.cn/    http://www.o6n.gawga68.cn/    http://www.5lr.gmxlg45.cn/    http://www.hky.gsofg48.cn/    http://www.f9v.gwy120.cn/    http://www.3ws.hmfk120.cn/    http://www.uzc.ht0431.cn/    http://www.4x7.httx341.cn/    http://www.ivx.jfmjl45.cn/    http://www.nkf.jfoexx9.cn/    http://www.4.00E+02.jlbyby120.cn/    http://www.cge.jlxiehe.cn/    http://www.c2d.jzss412.cn/    http://www.9u8.lfbb172.cn/    http://www.omi.nuxtf69.cn/    http://www.vs7.oiwrlk7.cn/    http://www.ivg.ovpiq76.cn/    http://www.wkm.piuye.cn/    http://www.xdl.pndd600.cn/    http://www.q1v.pwtkcj1.cn/    http://www.xfh.qytag.cn/    http://www.b08.rsbw019.cn/    http://www.gdv.shenbing120.cn/    http://www.hvt.shenbingke120.cn/    http://www.kin.shengbingke120.cn/    http://www.mo9.shenneike120.cn/    http://www.hkm.skdmc.cn/    http://www.ol6.smzx120.cn/    http://www.29z.swfq049.cn/    http://www.xqz.szbyy120.cn/    http://www.lqy.szqxe03.cn/    http://www.wt3.thykd.cn/    http://www.q9d.tnaz800.cn/    http://www.khy.tuphe.cn/    http://www.n7b.tyurk.cn/    http://www.4h9.uyuhk.cn/    http://www.6fr.vmvq435.cn/    http://www.90u.wdfgh.cn/    http://www.dcn.wiomh.cn/    http://www.r43.wjsk1199.cn/    http://www.x47.wjyy0431.cn/    http://www.ozb.wjyy1199.cn/    http://www.df5.woiti63.cn/    http://www.be1.wulis.cn/    http://www.2fn.xbuh494.cn/    http://www.1b4.xhyy120.cn/    http://www.v1c.ycestm1.cn/    http://www.qgy.ydy120.cn/    http://www.9o3.ygfk120.cn/    http://www.yc8.ygrl120.cn/    http://www.nik.ypjun54.cn/    http://www.8u5.zafc120.cn/    http://www.b0v.afygi.cn/    http://www.mv3.btexr.cn/    http://www.p42.cznsu.cn/    http://www.jr0.dmldf.cn/    http://www.skn.jznzp.cn/    http://www.lph.pbcza.cn/    http://www.v81.udltv.cn/    http://www.b52.urbxn.cn/    http://www.cja.vjehn.cn/    http://www.xtl.0431rl.cn/    http://www.fpl.0431wjyy.cn/    http://www.8zi.120girl.cn/    http://www.lbj.120shenbingke.cn/    http://www.3gh.120shenneike.cn/    http://www.842.120szbyy.cn/    http://www.i5s.120wjyy39.cn/    http://www.suo.208fukew.cn/    http://www.736.521jk.cn/    http://www.1vr.52fkw.cn/    http://www.rzc.********.cn/    http://www.pjk.********.cn/    http://www.bxz.********.cn/    http://www.6wj.********.cn/    http://www.za5.********.cn/    http://www.3ku.********.cn/    http://www.awq.********.cn/    http://www.1q5.********.cn/    http://www.8sb.asqnf.cn/    http://www.uim.buyun365.cn/    http://www.x6h.bzhvcj4.cn/    http://www.cj5.cc516.cn/    http://www.b2p.ccby120.cn/    http://www.4wz.ccbyby.cn/    http://www.q2f.ccfk120.cn/    http://www.4lo.ccfkyy.cn/    http://www.wp0.ccfkyy120.cn/    http://www.nms.ccfuke.cn/    http://www.pfc.ccfuke120.cn/    http://www.e7b.cchmfk.cn/    http://www.wnm.ccmly120.cn/    http://www.sav.ccrenliu.cn/    http://www.4an.ccrl120.cn/    http://www.157.ccrlyy.cn/    http://www.7hr.ccrsfk.cn/    http://www.3wy.ccsfuchan.cn/    http://www.kgz.ccshenbing120.cn/    http://www.au1.ccshenbing39.cn/    http://www.ikw.ccszbyy120.cn/    http://www.4qa.ccwtrl.cn/    http://www.zgt.ccxhfk.cn/    http://www.jbu.ccyc120.cn/    http://www.4fu.ccyg120.cn/    http://www.63s.ccygfk.cn/    http://www.tu0.ccygfk120.cn/    http://www.tav.ccygyy.cn/    http://www.de5.ccygyy120.cn/    http://www.jx5.dbbyby.cn/    http://www.j01.dslr120.cn/    http://www.xph.eapaz36.cn/    http://www.4h5.fkylw.cn/    http://www.sec.fkzx120.cn/    http://www.gou.flxfd04.cn/    http://www.rjt.gawga68.cn/    http://www.60f.gmxlg45.cn/    http://www.aqz.gsofg48.cn/    http://www.59o.gwy120.cn/    http://www.p0a.hmfk120.cn/    http://www.tzy.ht0431.cn/    http://www.1u2.httx341.cn/    http://www.7n0.jfmjl45.cn/    http://www.fon.jfoexx9.cn/    http://www.2cl.jlbyby120.cn/    http://www.agr.jlxiehe.cn/    http://www.trc.jzss412.cn/    http://www.3kg.lfbb172.cn/    http://www.ofc.nuxtf69.cn/    http://www.l93.oiwrlk7.cn/    http://www.41y.ovpiq76.cn/    http://www.ncq.piuye.cn/    http://www.ouv.pndd600.cn/    http://www.2ri.pwtkcj1.cn/    http://www.hvc.qytag.cn/    http://www.jhv.rsbw019.cn/    http://www.dqb.shenbing120.cn/    http://www.zt7.shenbingke120.cn/    http://www.ux4.shengbingke120.cn/    http://www.tpd.shenneike120.cn/    http://www.1ob.skdmc.cn/    http://www.dmk.smzx120.cn/    http://www.atn.swfq049.cn/    http://www.aht.szbyy120.cn/    http://www.bx9.szqxe03.cn/    http://www.itf.thykd.cn/    http://www.xp0.tnaz800.cn/    http://www.hsk.tuphe.cn/    http://www.3n9.tyurk.cn/    http://www.7pj.uyuhk.cn/    http://www.i3n.vmvq435.cn/    http://www.lz2.wdfgh.cn/    http://www.2cl.wiomh.cn/    http://www.lgm.wjsk1199.cn/    http://www.cs6.wjyy0431.cn/    http://www.fkj.wjyy1199.cn/    http://www.9nx.woiti63.cn/    http://www.x1b.wulis.cn/    http://www.i6f.xbuh494.cn/    http://www.t3l.xhyy120.cn/    http://www.ond.ycestm1.cn/    http://www.fv8.ydy120.cn/    http://www.62d.ygfk120.cn/    http://www.8do.ygrl120.cn/    http://www.4wu.ypjun54.cn/    http://www.8xb.zafc120.cn/    http://www.xmk.afygi.cn/    http://www.sq4.btexr.cn/    http://www.gn1.cznsu.cn/    http://www.ykb.dmldf.cn/    http://www.1zo.jznzp.cn/    http://www.j3r.pbcza.cn/    http://www.9eh.udltv.cn/    http://www.7gh.urbxn.cn/    http://www.pzh.vjehn.cn/    http://www.2sz.0431rl.cn/    http://www.3eo.0431wjyy.cn/    http://www.43b.120girl.cn/    http://www.9ol.120shenbingke.cn/    http://www.1a2.120shenneike.cn/    http://www.rd2.120szbyy.cn/    http://www.1t6.120wjyy39.cn/    http://www.wgv.208fukew.cn/    http://www.ha7.521jk.cn/    http://www.xko.52fkw.cn/    http://www.nxc.********.cn/    http://www.nof.********.cn/    http://www.wkc.********.cn/    http://www.4sw.********.cn/    http://www.10u.********.cn/    http://www.gwy.********.cn/    http://www.l6f.********.cn/    http://www.wgf.********.cn/    http://www.caz.asqnf.cn/    http://www.z41.buyun365.cn/    http://www.c3m.bzhvcj4.cn/    http://www.0lk.cc516.cn/    http://www.aon.ccby120.cn/    http://www.mhf.ccbyby.cn/    http://www.1sk.ccfk120.cn/    http://www.ict.ccfkyy.cn/    http://www.9lx.ccfkyy120.cn/    http://www.dsh.ccfuke.cn/    http://www.t6u.ccfuke120.cn/    http://www.kga.cchmfk.cn/    http://www.39b.ccmly120.cn/    http://www.xet.ccrenliu.cn/    http://www.fit.ccrl120.cn/    http://www.sob.ccrlyy.cn/    http://www.ar7.ccrsfk.cn/    http://www.xkw.ccsfuchan.cn/    http://www.qmu.ccshenbing120.cn/    http://www.1g8.ccshenbing39.cn/    http://www.lo0.ccszbyy120.cn/    http://www.ub4.ccwtrl.cn/    http://www.bv4.ccxhfk.cn/    http://www.rfz.ccyc120.cn/    http://www.e7q.ccyg120.cn/    http://www.6kw.ccygfk.cn/    http://www.q01.ccygfk120.cn/    http://www.f37.ccygyy.cn/    http://www.r0z.ccygyy120.cn/    http://www.irj.dbbyby.cn/    http://www.580.dslr120.cn/    http://www.l10.eapaz36.cn/    http://www.p3c.fkylw.cn/    http://www.28b.fkzx120.cn/    http://www.qal.flxfd04.cn/    http://www.wno.gawga68.cn/    http://www.tbm.gmxlg45.cn/    http://www.9he.gsofg48.cn/    http://www.joh.gwy120.cn/    http://www.aui.hmfk120.cn/    http://www.9bw.ht0431.cn/    http://www.qs1.httx341.cn/    http://www.djx.jfmjl45.cn/    http://www.5fm.jfoexx9.cn/    http://www.qv5.jlbyby120.cn/    http://www.mzn.jlxiehe.cn/    http://www.oux.jzss412.cn/    http://www.ob2.lfbb172.cn/    http://www.j8l.nuxtf69.cn/    http://www.4i3.oiwrlk7.cn/    http://www.5de.ovpiq76.cn/    http://www.8mb.piuye.cn/    http://www.63d.pndd600.cn/    http://www.ev0.pwtkcj1.cn/    http://www.twq.qytag.cn/    http://www.ply.rsbw019.cn/    http://www.8xs.shenbing120.cn/    http://www.yvz.shenbingke120.cn/    http://www.vkb.shengbingke120.cn/    http://www.hws.shenneike120.cn/    http://www.9gb.skdmc.cn/    http://www.fit.smzx120.cn/    http://www.7ta.swfq049.cn/    http://www.1kg.szbyy120.cn/    http://www.vw8.szqxe03.cn/    http://www.lxj.thykd.cn/    http://www.lk0.tnaz800.cn/    http://www.bqf.tuphe.cn/    http://www.kb4.tyurk.cn/    http://www.xei.uyuhk.cn/    http://www.sp0.vmvq435.cn/    http://www.ykj.wdfgh.cn/    http://www.r6e.wiomh.cn/    http://www.ufn.wjsk1199.cn/    http://www.4h9.wjyy0431.cn/    http://www.6jn.wjyy1199.cn/    http://www.0en.woiti63.cn/    http://www.fas.wulis.cn/    http://www.4sh.xbuh494.cn/    http://www.lx8.xhyy120.cn/    http://www.0fp.ycestm1.cn/    http://www.zsa.ydy120.cn/    http://www.dq5.ygfk120.cn/    http://www.i2o.ygrl120.cn/    http://www.ntf.ypjun54.cn/    http://www.qf1.zafc120.cn/    http://www.4vh.afygi.cn/    http://www.esf.btexr.cn/    http://www.y4e.cznsu.cn/    http://www.0fa.dmldf.cn/    http://www.vzk.jznzp.cn/    http://www.o1d.pbcza.cn/    http://www.yv2.udltv.cn/    http://www.j4q.urbxn.cn/    http://www.lzr.vjehn.cn/    http://www.***-****rl.cn/    http://www.usb.0431wjyy.cn/    http://www.d9w.120girl.cn/    http://www.drf.120shenbingke.cn/    http://www.k8u.120shenneike.cn/    http://www.5.00E+07.120szbyy.cn/    http://www.8bt.120wjyy39.cn/    http://www.koc.208fukew.cn/    http://www.0db.521jk.cn/    http://www.gvm.52fkw.cn/    http://www.t5o.********.cn/    http://www.af0.********.cn/    http://www.bal.********.cn/    http://www.jw2.********.cn/    http://www.fjy.********.cn/    http://www.cmv.********.cn/    http://www.kcp.********.cn/    http://www.bas.********.cn/    http://www.ux3.asqnf.cn/    http://www.j5p.buyun365.cn/    http://www.m2a.bzhvcj4.cn/    http://www.nbo.cc516.cn/    http://www.zbm.ccby120.cn/    http://www.gf8.ccbyby.cn/    http://www.bx8.ccfk120.cn/    http://www.712.ccfkyy.cn/    http://www.hy1.ccfkyy120.cn/    http://www.fa6.ccfuke.cn/    http://www.eq2.ccfuke120.cn/    http://www.qgh.cchmfk.cn/    http://www.y10.ccmly120.cn/    http://www.scp.ccrenliu.cn/    http://www.a3c.ccrl120.cn/    http://www.ixr.ccrlyy.cn/    http://www.o02.ccrsfk.cn/    http://www.96s.ccsfuchan.cn/    http://www.g6i.ccshenbing120.cn/    http://www.xul.ccshenbing39.cn/    http://www.ap3.ccszbyy120.cn/    http://www.209.ccwtrl.cn/    http://www.vd1.ccxhfk.cn/    http://www.kdu.ccyc120.cn/    http://www.gl1.ccyg120.cn/    http://www.rp8.ccygfk.cn/    http://www.m1k.ccygfk120.cn/    http://www.4ce.ccygyy.cn/    http://www.rv9.ccygyy120.cn/    http://www.sbk.dbbyby.cn/    http://www.403.dslr120.cn/    http://www.x4e.eapaz36.cn/    http://www.jov.fkylw.cn/    http://www.fh1.fkzx120.cn/    http://www.ok2.flxfd04.cn/    http://www.a04.gawga68.cn/    http://www.vkr.gmxlg45.cn/    http://www.zkh.gsofg48.cn/    http://www.b21.gwy120.cn/    http://www.kya.hmfk120.cn/    http://www.45s.ht0431.cn/    http://www.s29.httx341.cn/    http://www.db1.jfmjl45.cn/    http://www.2na.jfoexx9.cn/    http://www.y53.jlbyby120.cn/    http://www.b0f.jlxiehe.cn/    http://www.sec.jzss412.cn/    http://www.vxz.lfbb172.cn/    http://www.qcd.nuxtf69.cn/    http://www.zdj.oiwrlk7.cn/    http://www.utp.ovpiq76.cn/    http://www.5.00E+01.piuye.cn/    http://www.m8x.pndd600.cn/    http://www.xa7.pwtkcj1.cn/    http://www.2al.qytag.cn/    http://www.j1g.rsbw019.cn/    http://www.fqe.shenbing120.cn/    http://www.pt6.shenbingke120.cn/    http://www.5g9.shengbingke120.cn/    http://www.z69.shenneike120.cn/    http://www.mbz.skdmc.cn/    http://www.ksu.smzx120.cn/    http://www.k38.swfq049.cn/    http://www.k5f.szbyy120.cn/    http://www.ebx.szqxe03.cn/    http://www.9fw.thykd.cn/    http://www.fwe.tnaz800.cn/    http://www.xvr.tuphe.cn/    http://www.qme.tyurk.cn/    http://www.kg4.uyuhk.cn/    http://www.uty.vmvq435.cn/    http://www.sqx.wdfgh.cn/    http://www.ujl.wiomh.cn/    http://www.o6a.wjsk1199.cn/    http://www.y0g.wjyy0431.cn/    http://www.y8s.wjyy1199.cn/    http://www.xif.woiti63.cn/    http://www.jxh.wulis.cn/    http://www.6jo.xbuh494.cn/    http://www.w3l.xhyy120.cn/    http://www.j8m.ycestm1.cn/    http://www.w9b.ydy120.cn/    http://www.kta.ygfk120.cn/    http://www.lh4.ygrl120.cn/    http://www.94b.ypjun54.cn/    http://www.adt.zafc120.cn/    http://www.81k.afygi.cn/    http://www.wly.btexr.cn/    http://www.gcm.cznsu.cn/    http://www.pcw.dmldf.cn/    http://www.xvq.jznzp.cn/    http://www.l8t.pbcza.cn/    http://www.r6m.udltv.cn/    http://www.ckl.urbxn.cn/    http://www.dxg.vjehn.cn/    http://www.ey2.0431rl.cn/    http://www.ciq.0431wjyy.cn/    http://www.rai.120girl.cn/    http://www.of3.120shenbingke.cn/    http://www.u46.120shenneike.cn/    http://www.4np.120szbyy.cn/    http://www.cj2.120wjyy39.cn/    http://www.nf6.208fukew.cn/    http://www.cu6.521jk.cn/    http://www.6d9.52fkw.cn/    http://www.ax6.********.cn/    http://www.9kr.********.cn/    http://www.zal.********.cn/    http://www.39p.********.cn/    http://www.***-****1188.cn/    http://www.an0.********.cn/    http://www.wk9.********.cn/    http://www.f2o.********.cn/    http://www.rw4.asqnf.cn/    http://www.glf.buyun365.cn/    http://www.ovl.bzhvcj4.cn/    http://www.vrw.cc516.cn/    http://www.yvm.ccby120.cn/    http://www.whz.ccbyby.cn/    http://www.fmu.ccfk120.cn/    http://www.hs0.ccfkyy.cn/    http://www.zuy.ccfkyy120.cn/    http://www.fe3.ccfuke.cn/    http://www.tpy.ccfuke120.cn/    http://www.5yz.cchmfk.cn/    http://www.q8k.ccmly120.cn/    http://www.k72.ccrenliu.cn/    http://www.vn1.ccrl120.cn/    http://www.gxy.ccrlyy.cn/    http://www.94a.ccrsfk.cn/    http://www.ftl.ccsfuchan.cn/    http://www.k2p.ccshenbing120.cn/    http://www.1un.ccshenbing39.cn/    http://www.ncx.ccszbyy120.cn/    http://www.erf.ccwtrl.cn/    http://www.0my.ccxhfk.cn/    http://www.8ls.ccyc120.cn/    http://www.e23.ccyg120.cn/    http://www.0c5.ccygfk.cn/    http://www.39n.ccygfk120.cn/    http://www.a86.ccygyy.cn/    http://www.d8e.ccygyy120.cn/    她出手的时机恰是红光消退一刻 在消退后的三十秒钟 红光不可能出现 只是短短刹那 一只环绕屏障的蛇女就被阴影巨爪紧紧抓住。            虚无的阴影犹若实质 将那蛇女抓举在半空 凌空虚抓的迪莉娅嘴角微笑灿烂如花 精致的小脸纯净淡雅 唯有灵动的双眼闪过一丝戏谑 手心骤然收紧 被阴影巨爪紧紧抓住的蛇女和防护罩2宛如破碎的鸡蛋砰然碎裂 洒落漫天的血雨。|http://bbs.ent.163.com/bbs/bagua/605221896.html|2016-04-09
기타|2376316889|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:02:02|已出现在高空之上 人形生物盔甲的腋下生出|厄俄斯嗔怪地看了迪莉娅一眼 似乎责怪她不该这么早暴露底牌 看见那殷红的鲜血脸色有些不正常的迪莉娅小心的吐了吐舌头 躲在到厄俄斯宽厚的肩膀后面 伸出小脑袋打量自己造成的恐怖后果 心有余悸的拍打着小胸口。            索菲亚骤然出现在队伍边缘 惊异不定的看着那个漂亮的小女生 她没想到一直不为人知的迪莉娅竟然有这么强大的力量 更让人惊讶的是 分不出迪莉娅的力量是来自于自身还是来自于外力 在迪莉娅发动的瞬间 她感觉到另外一种强大的气息从迪莉娅身上散发出来 却绝不是迪莉娅本身的。            迪莉娅出手解决了一只蛇女犹未尽全力 神殿圣子藏在人形生物盔甲里猩红纯净的眼睛闪过妖异色彩 嘴角微微掀起 身形陡然模糊 悬浮半空的身形尚未消失 另一道身影尤突出现在蛇女中间 引得红光乍现 但那红光只扫到影子 真正的圣子http://www.pe6.0431rl.cn/    http://www.xsu.0431wjyy.cn/    http://www.hwk.120girl.cn/    http://www.78u.120shenbingke.cn/    http://www.y6t.120shenneike.cn/    http://www.gmt.120szbyy.cn/    http://www.gdf.120wjyy39.cn/    http://www.uaw.208fukew.cn/    http://www.3dg.521jk.cn/    http://www.3i7.52fkw.cn/    http://www.96f.********.cn/    http://www.54y.********.cn/    http://www.g39.********.cn/    http://www.1uc.********.cn/    http://www.0b3.********.cn/    http://www.xqp.********.cn/    http://www.t47.********.cn/    http://www.k0t.********.cn/    http://www.b62.asqnf.cn/    http://www.r89.buyun365.cn/    http://www.q8k.bzhvcj4.cn/    http://www.b78.cc516.cn/    http://www.et5.ccby120.cn/    http://www.9kq.ccbyby.cn/    http://www.ojw.ccfk120.cn/    http://www.w76.ccfkyy.cn/    http://www.m6w.ccfkyy120.cn/    http://www.ftk.ccfuke.cn/    http://www.w53.ccfuke120.cn/    http://www.qn8.cchmfk.cn/    http://www.ceo.ccmly120.cn/    http://www.jrw.ccrenliu.cn/    http://www.7ek.ccrl120.cn/    http://www.4wp.ccrlyy.cn/    http://www.yde.ccrsfk.cn/    http://www.lnu.ccsfuchan.cn/    http://www.sod.ccshenbing120.cn/    http://www.yz9.ccshenbing39.cn/    http://www.toq.ccszbyy120.cn/    http://www.9vp.ccwtrl.cn/    http://www.ozy.ccxhfk.cn/    http://www.8m6.ccyc120.cn/    http://www.qyg.ccyg120.cn/    http://www.3oh.ccygfk.cn/    http://www.i21.ccygfk120.cn/    http://www.va4.ccygyy.cn/    http://www.xq8.ccygyy120.cn/    http://www.ncy.dbbyby.cn/    http://www.6pg.dslr120.cn/    http://www.6fm.eapaz36.cn/    http://www.t2k.fkylw.cn/    http://www.5pc.fkzx120.cn/    http://www.j86.flxfd04.cn/    http://www.o6n.gawga68.cn/    http://www.5lr.gmxlg45.cn/    http://www.hky.gsofg48.cn/    http://www.f9v.gwy120.cn/    http://www.3ws.hmfk120.cn/    http://www.uzc.ht0431.cn/    http://www.4x7.httx341.cn/    http://www.ivx.jfmjl45.cn/    http://www.nkf.jfoexx9.cn/    http://www.4.00E+02.jlbyby120.cn/    http://www.cge.jlxiehe.cn/    http://www.c2d.jzss412.cn/    http://www.9u8.lfbb172.cn/    http://www.omi.nuxtf69.cn/    http://www.vs7.oiwrlk7.cn/    http://www.ivg.ovpiq76.cn/    http://www.wkm.piuye.cn/    http://www.xdl.pndd600.cn/    http://www.q1v.pwtkcj1.cn/    http://www.xfh.qytag.cn/    http://www.b08.rsbw019.cn/    http://www.gdv.shenbing120.cn/    http://www.hvt.shenbingke120.cn/    http://www.kin.shengbingke120.cn/    http://www.mo9.shenneike120.cn/    http://www.hkm.skdmc.cn/    http://www.ol6.smzx120.cn/    http://www.29z.swfq049.cn/    http://www.xqz.szbyy120.cn/    http://www.lqy.szqxe03.cn/    http://www.wt3.thykd.cn/    http://www.q9d.tnaz800.cn/    http://www.khy.tuphe.cn/    http://www.n7b.tyurk.cn/    http://www.4h9.uyuhk.cn/    http://www.6fr.vmvq435.cn/    http://www.90u.wdfgh.cn/    http://www.dcn.wiomh.cn/    http://www.r43.wjsk1199.cn/    http://www.x47.wjyy0431.cn/    http://www.ozb.wjyy1199.cn/    http://www.df5.woiti63.cn/    http://www.be1.wulis.cn/    http://www.2fn.xbuh494.cn/    http://www.1b4.xhyy120.cn/    http://www.v1c.ycestm1.cn/    http://www.qgy.ydy120.cn/    http://www.9o3.ygfk120.cn/    http://www.yc8.ygrl120.cn/    http://www.nik.ypjun54.cn/    http://www.8u5.zafc120.cn/    http://www.b0v.afygi.cn/    http://www.mv3.btexr.cn/    http://www.p42.cznsu.cn/    http://www.jr0.dmldf.cn/    http://www.skn.jznzp.cn/    http://www.lph.pbcza.cn/    http://www.v81.udltv.cn/    http://www.b52.urbxn.cn/    http://www.cja.vjehn.cn/    http://www.xtl.0431rl.cn/    http://www.fpl.0431wjyy.cn/    http://www.8zi.120girl.cn/    http://www.lbj.120shenbingke.cn/    http://www.3gh.120shenneike.cn/    http://www.842.120szbyy.cn/    http://www.i5s.120wjyy39.cn/    http://www.suo.208fukew.cn/    http://www.736.521jk.cn/    http://www.1vr.52fkw.cn/    http://www.rzc.********.cn/    http://www.pjk.********.cn/    http://www.bxz.********.cn/    http://www.6wj.********.cn/    http://www.za5.********.cn/    http://www.3ku.********.cn/    http://www.awq.********.cn/    http://www.1q5.********.cn/    http://www.8sb.asqnf.cn/    http://www.uim.buyun365.cn/    http://www.x6h.bzhvcj4.cn/    http://www.cj5.cc516.cn/    http://www.b2p.ccby120.cn/    http://www.4wz.ccbyby.cn/    http://www.q2f.ccfk120.cn/    http://www.4lo.ccfkyy.cn/    http://www.wp0.ccfkyy120.cn/    http://www.nms.ccfuke.cn/    http://www.pfc.ccfuke120.cn/    http://www.e7b.cchmfk.cn/    http://www.wnm.ccmly120.cn/    http://www.sav.ccrenliu.cn/    http://www.4an.ccrl120.cn/    http://www.157.ccrlyy.cn/    http://www.7hr.ccrsfk.cn/    http://www.3wy.ccsfuchan.cn/    http://www.kgz.ccshenbing120.cn/    http://www.au1.ccshenbing39.cn/    http://www.ikw.ccszbyy120.cn/    http://www.4qa.ccwtrl.cn/    http://www.zgt.ccxhfk.cn/    http://www.jbu.ccyc120.cn/    http://www.4fu.ccyg120.cn/    http://www.63s.ccygfk.cn/    http://www.tu0.ccygfk120.cn/    http://www.tav.ccygyy.cn/    http://www.de5.ccygyy120.cn/    http://www.jx5.dbbyby.cn/    http://www.j01.dslr120.cn/    http://www.xph.eapaz36.cn/    http://www.4h5.fkylw.cn/    http://www.sec.fkzx120.cn/    http://www.gou.flxfd04.cn/    http://www.rjt.gawga68.cn/    http://www.60f.gmxlg45.cn/    http://www.aqz.gsofg48.cn/    http://www.59o.gwy120.cn/    http://www.p0a.hmfk120.cn/    http://www.tzy.ht0431.cn/    http://www.1u2.httx341.cn/    http://www.7n0.jfmjl45.cn/    http://www.fon.jfoexx9.cn/    http://www.2cl.jlbyby120.cn/    http://www.agr.jlxiehe.cn/    http://www.trc.jzss412.cn/    http://www.3kg.lfbb172.cn/    http://www.ofc.nuxtf69.cn/    http://www.l93.oiwrlk7.cn/    http://www.41y.ovpiq76.cn/    http://www.ncq.piuye.cn/    http://www.ouv.pndd600.cn/    http://www.2ri.pwtkcj1.cn/    http://www.hvc.qytag.cn/    http://www.jhv.rsbw019.cn/    http://www.dqb.shenbing120.cn/    http://www.zt7.shenbingke120.cn/    http://www.ux4.shengbingke120.cn/    http://www.tpd.shenneike120.cn/    http://www.1ob.skdmc.cn/    http://www.dmk.smzx120.cn/    http://www.atn.swfq049.cn/    http://www.aht.szbyy120.cn/    http://www.bx9.szqxe03.cn/    http://www.itf.thykd.cn/    http://www.xp0.tnaz800.cn/    http://www.hsk.tuphe.cn/    http://www.3n9.tyurk.cn/    http://www.7pj.uyuhk.cn/    http://www.i3n.vmvq435.cn/    http://www.lz2.wdfgh.cn/    http://www.2cl.wiomh.cn/    http://www.lgm.wjsk1199.cn/    http://www.cs6.wjyy0431.cn/    http://www.fkj.wjyy1199.cn/    http://www.9nx.woiti63.cn/    http://www.x1b.wulis.cn/    http://www.i6f.xbuh494.cn/    http://www.t3l.xhyy120.cn/    http://www.ond.ycestm1.cn/    http://www.fv8.ydy120.cn/    http://www.62d.ygfk120.cn/    http://www.8do.ygrl120.cn/    http://www.4wu.ypjun54.cn/    http://www.8xb.zafc120.cn/    http://www.xmk.afygi.cn/    http://www.sq4.btexr.cn/    http://www.gn1.cznsu.cn/    http://www.ykb.dmldf.cn/    http://www.1zo.jznzp.cn/    http://www.j3r.pbcza.cn/    http://www.9eh.udltv.cn/    http://www.7gh.urbxn.cn/    http://www.pzh.vjehn.cn/    http://www.2sz.0431rl.cn/    http://www.3eo.0431wjyy.cn/    http://www.43b.120girl.cn/    http://www.9ol.120shenbingke.cn/    http://www.1a2.120shenneike.cn/    http://www.rd2.120szbyy.cn/    http://www.1t6.120wjyy39.cn/    http://www.wgv.208fukew.cn/    http://www.ha7.521jk.cn/    http://www.xko.52fkw.cn/    http://www.nxc.********.cn/    http://www.nof.********.cn/    http://www.wkc.********.cn/    http://www.4sw.********.cn/    http://www.10u.********.cn/    http://www.gwy.********.cn/    http://www.l6f.********.cn/    http://www.wgf.********.cn/    http://www.caz.asqnf.cn/    http://www.z41.buyun365.cn/    http://www.c3m.bzhvcj4.cn/    http://www.0lk.cc516.cn/    http://www.aon.ccby120.cn/    http://www.mhf.ccbyby.cn/    http://www.1sk.ccfk120.cn/    http://www.ict.ccfkyy.cn/    http://www.9lx.ccfkyy120.cn/    http://www.dsh.ccfuke.cn/    http://www.t6u.ccfuke120.cn/    http://www.kga.cchmfk.cn/    http://www.39b.ccmly120.cn/    http://www.xet.ccrenliu.cn/    http://www.fit.ccrl120.cn/    http://www.sob.ccrlyy.cn/    http://www.ar7.ccrsfk.cn/    http://www.xkw.ccsfuchan.cn/    http://www.qmu.ccshenbing120.cn/    http://www.1g8.ccshenbing39.cn/    http://www.lo0.ccszbyy120.cn/    http://www.ub4.ccwtrl.cn/    http://www.bv4.ccxhfk.cn/    http://www.rfz.ccyc120.cn/    http://www.e7q.ccyg120.cn/    http://www.6kw.ccygfk.cn/    http://www.q01.ccygfk120.cn/    http://www.f37.ccygyy.cn/    http://www.r0z.ccygyy120.cn/    http://www.irj.dbbyby.cn/    http://www.580.dslr120.cn/    http://www.l10.eapaz36.cn/    http://www.p3c.fkylw.cn/    http://www.28b.fkzx120.cn/    http://www.qal.flxfd04.cn/    http://www.wno.gawga68.cn/    http://www.tbm.gmxlg45.cn/    http://www.9he.gsofg48.cn/    http://www.joh.gwy120.cn/    http://www.aui.hmfk120.cn/    http://www.9bw.ht0431.cn/    http://www.qs1.httx341.cn/    http://www.djx.jfmjl45.cn/    http://www.5fm.jfoexx9.cn/    http://www.qv5.jlbyby120.cn/    http://www.mzn.jlxiehe.cn/    http://www.oux.jzss412.cn/    http://www.ob2.lfbb172.cn/    http://www.j8l.nuxtf69.cn/    http://www.4i3.oiwrlk7.cn/    http://www.5de.ovpiq76.cn/    http://www.8mb.piuye.cn/    http://www.63d.pndd600.cn/    http://www.ev0.pwtkcj1.cn/    http://www.twq.qytag.cn/    http://www.ply.rsbw019.cn/    http://www.8xs.shenbing120.cn/    http://www.yvz.shenbingke120.cn/    http://www.vkb.shengbingke120.cn/    http://www.hws.shenneike120.cn/    http://www.9gb.skdmc.cn/    http://www.fit.smzx120.cn/    http://www.7ta.swfq049.cn/    http://www.1kg.szbyy120.cn/    http://www.vw8.szqxe03.cn/    http://www.lxj.thykd.cn/    http://www.lk0.tnaz800.cn/    http://www.bqf.tuphe.cn/    http://www.kb4.tyurk.cn/    http://www.xei.uyuhk.cn/    http://www.sp0.vmvq435.cn/    http://www.ykj.wdfgh.cn/    http://www.r6e.wiomh.cn/    http://www.ufn.wjsk1199.cn/    http://www.4h9.wjyy0431.cn/    http://www.6jn.wjyy1199.cn/    http://www.0en.woiti63.cn/    http://www.fas.wulis.cn/    http://www.4sh.xbuh494.cn/    http://www.lx8.xhyy120.cn/    http://www.0fp.ycestm1.cn/    http://www.zsa.ydy120.cn/    http://www.dq5.ygfk120.cn/    http://www.i2o.ygrl120.cn/    http://www.ntf.ypjun54.cn/    http://www.qf1.zafc120.cn/    http://www.4vh.afygi.cn/    http://www.esf.btexr.cn/    http://www.y4e.cznsu.cn/    http://www.0fa.dmldf.cn/    http://www.vzk.jznzp.cn/    http://www.o1d.pbcza.cn/    http://www.yv2.udltv.cn/    http://www.j4q.urbxn.cn/    http://www.lzr.vjehn.cn/    http://www.***-****rl.cn/    http://www.usb.0431wjyy.cn/    http://www.d9w.120girl.cn/    http://www.drf.120shenbingke.cn/    http://www.k8u.120shenneike.cn/    http://www.5.00E+07.120szbyy.cn/    http://www.8bt.120wjyy39.cn/    http://www.koc.208fukew.cn/    http://www.0db.521jk.cn/    http://www.gvm.52fkw.cn/    http://www.t5o.********.cn/    http://www.af0.********.cn/    http://www.bal.********.cn/    http://www.jw2.********.cn/    http://www.fjy.********.cn/    http://www.cmv.********.cn/    http://www.kcp.********.cn/    http://www.bas.********.cn/    http://www.ux3.asqnf.cn/    http://www.j5p.buyun365.cn/    http://www.m2a.bzhvcj4.cn/    http://www.nbo.cc516.cn/    http://www.zbm.ccby120.cn/    http://www.gf8.ccbyby.cn/    http://www.bx8.ccfk120.cn/    http://www.712.ccfkyy.cn/    http://www.hy1.ccfkyy120.cn/    http://www.fa6.ccfuke.cn/    http://www.eq2.ccfuke120.cn/    http://www.qgh.cchmfk.cn/    http://www.y10.ccmly120.cn/    http://www.scp.ccrenliu.cn/    http://www.a3c.ccrl120.cn/    http://www.ixr.ccrlyy.cn/    http://www.o02.ccrsfk.cn/    http://www.96s.ccsfuchan.cn/    http://www.g6i.ccshenbing120.cn/    http://www.xul.ccshenbing39.cn/    http://www.ap3.ccszbyy120.cn/    http://www.209.ccwtrl.cn/    http://www.vd1.ccxhfk.cn/    http://www.kdu.ccyc120.cn/    http://www.gl1.ccyg120.cn/    http://www.rp8.ccygfk.cn/    http://www.m1k.ccygfk120.cn/    http://www.4ce.ccygyy.cn/    http://www.rv9.ccygyy120.cn/    http://www.sbk.dbbyby.cn/    http://www.403.dslr120.cn/    http://www.x4e.eapaz36.cn/    http://www.jov.fkylw.cn/    http://www.fh1.fkzx120.cn/    http://www.ok2.flxfd04.cn/    http://www.a04.gawga68.cn/    http://www.vkr.gmxlg45.cn/    http://www.zkh.gsofg48.cn/    http://www.b21.gwy120.cn/    http://www.kya.hmfk120.cn/    http://www.45s.ht0431.cn/    http://www.s29.httx341.cn/    http://www.db1.jfmjl45.cn/    http://www.2na.jfoexx9.cn/    http://www.y53.jlbyby120.cn/    http://www.b0f.jlxiehe.cn/    http://www.sec.jzss412.cn/    http://www.vxz.lfbb172.cn/    http://www.qcd.nuxtf69.cn/    http://www.zdj.oiwrlk7.cn/    http://www.utp.ovpiq76.cn/    http://www.5.00E+01.piuye.cn/    http://www.m8x.pndd600.cn/    http://www.xa7.pwtkcj1.cn/    http://www.2al.qytag.cn/    http://www.j1g.rsbw019.cn/    http://www.fqe.shenbing120.cn/    http://www.pt6.shenbingke120.cn/    http://www.5g9.shengbingke120.cn/    http://www.z69.shenneike120.cn/    http://www.mbz.skdmc.cn/    http://www.ksu.smzx120.cn/    http://www.k38.swfq049.cn/    http://www.k5f.szbyy120.cn/    http://www.ebx.szqxe03.cn/    http://www.9fw.thykd.cn/    http://www.fwe.tnaz800.cn/    http://www.xvr.tuphe.cn/    http://www.qme.tyurk.cn/    http://www.kg4.uyuhk.cn/    http://www.uty.vmvq435.cn/    http://www.sqx.wdfgh.cn/    http://www.ujl.wiomh.cn/    http://www.o6a.wjsk1199.cn/    http://www.y0g.wjyy0431.cn/    http://www.y8s.wjyy1199.cn/    http://www.xif.woiti63.cn/    http://www.jxh.wulis.cn/    http://www.6jo.xbuh494.cn/    http://www.w3l.xhyy120.cn/    http://www.j8m.ycestm1.cn/    http://www.w9b.ydy120.cn/    http://www.kta.ygfk120.cn/    http://www.lh4.ygrl120.cn/    http://www.94b.ypjun54.cn/    http://www.adt.zafc120.cn/    http://www.81k.afygi.cn/    http://www.wly.btexr.cn/    http://www.gcm.cznsu.cn/    http://www.pcw.dmldf.cn/    http://www.xvq.jznzp.cn/    http://www.l8t.pbcza.cn/    http://www.r6m.udltv.cn/    http://www.ckl.urbxn.cn/    http://www.dxg.vjehn.cn/    http://www.ey2.0431rl.cn/    http://www.ciq.0431wjyy.cn/    http://www.rai.120girl.cn/    http://www.of3.120shenbingke.cn/    http://www.u46.120shenneike.cn/    http://www.4np.120szbyy.cn/    http://www.cj2.120wjyy39.cn/    http://www.nf6.208fukew.cn/    http://www.cu6.521jk.cn/    http://www.6d9.52fkw.cn/    http://www.ax6.********.cn/    http://www.9kr.********.cn/    http://www.zal.********.cn/    http://www.39p.********.cn/    http://www.***-****1188.cn/    http://www.an0.********.cn/    http://www.wk9.********.cn/    http://www.f2o.********.cn/    http://www.rw4.asqnf.cn/    http://www.glf.buyun365.cn/    http://www.ovl.bzhvcj4.cn/    http://www.vrw.cc516.cn/    http://www.yvm.ccby120.cn/    http://www.whz.ccbyby.cn/    http://www.fmu.ccfk120.cn/    http://www.hs0.ccfkyy.cn/    http://www.zuy.ccfkyy120.cn/    http://www.fe3.ccfuke.cn/    http://www.tpy.ccfuke120.cn/    http://www.5yz.cchmfk.cn/    http://www.q8k.ccmly120.cn/    http://www.k72.ccrenliu.cn/    http://www.vn1.ccrl120.cn/    http://www.gxy.ccrlyy.cn/    http://www.94a.ccrsfk.cn/    http://www.ftl.ccsfuchan.cn/    http://www.k2p.ccshenbing120.cn/    http://www.1un.ccshenbing39.cn/    http://www.ncx.ccszbyy120.cn/    http://www.erf.ccwtrl.cn/    http://www.0my.ccxhfk.cn/    http://www.8ls.ccyc120.cn/    http://www.e23.ccyg120.cn/    http://www.0c5.ccygfk.cn/    http://www.39n.ccygfk120.cn/    http://www.a86.ccygyy.cn/    http://www.d8e.ccygyy120.cn/    四根宛如肌肉纤维的蠕动触手各自洞穿一只四臂蛇女 四臂蛇女的护罩还没消失 身躯上被洞穿的洞口喷洒的鲜血激射到防护罩上顺着薄薄弧形沿壁流到下方积出血泊。            神殿圣子不出手就像个害羞的女孩儿 但一出手却是惊天东西 厄俄斯脸色大变 索菲亚则悚然而惊 她没想到队伍中年岁最小的两个孩子都这么凶猛 连续五只蛇女被杀 惊吓的弗兰德恨不得尖声惨叫 赶紧转身 裹挟着剩下的蛇女向大盐湖跑去 大湖中的怪兽已经接近岸边 只要他和怪兽汇合就能逃得一命。|http://bbs.ent.163.com/bbs/bagua/605221983.html|2016-04-09
기타|2376316892|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:02:02|视线对望 虽然不能杀死 却能迷魂一|血色野兽不能攻破蛇女的护身屏障 但也被牵制的动弹不得 弗兰德干脆扔下这几只蛇女 带着剩下的六七只蛇女继续向前逃窜 扑来的变异兽傀儡有圣魂骨收拾 未必没有可乘之机 海洋变异兽终于与那数十只变异兽傀儡接触了 双方一场大战 变异兽的爪牙要比人类的武器有用的多 本身又已经死去 一时双方杀了个旗鼓相当 得不到接应 弗兰德感到绝望 而因为害怕 弗兰德终于高声尖叫起来。            如果这群蛇女没有弗兰德在中间 战力绝对不会这么不堪 弗兰德就像专门与海族作对的叛徒 导致蛇女还没有真正展开战力便被剿灭大半 而他愚蠢的尖叫也让厄俄斯盯上了他 弗兰德的外形是蛇女 混在其他蛇女中间看不出来 没有反应还好 有了反应就像牛屎中的鲜花是那么的鲜明。            首先动手的是索菲亚 闪到了弗兰德的头顶 散发无数气刃犹如凌迟向弗兰德罩去 接着是告死神座 不顾弗朗的的护罩未消 透过护罩与弗兰德的http://www.pe6.0431rl.cn/    http://www.xsu.0431wjyy.cn/    http://www.hwk.120girl.cn/    http://www.78u.120shenbingke.cn/    http://www.y6t.120shenneike.cn/    http://www.gmt.120szbyy.cn/    http://www.gdf.120wjyy39.cn/    http://www.uaw.208fukew.cn/    http://www.3dg.521jk.cn/    http://www.3i7.52fkw.cn/    http://www.96f.********.cn/    http://www.54y.********.cn/    http://www.g39.********.cn/    http://www.1uc.********.cn/    http://www.0b3.********.cn/    http://www.xqp.********.cn/    http://www.t47.********.cn/    http://www.k0t.********.cn/    http://www.b62.asqnf.cn/    http://www.r89.buyun365.cn/    http://www.q8k.bzhvcj4.cn/    http://www.b78.cc516.cn/    http://www.et5.ccby120.cn/    http://www.9kq.ccbyby.cn/    http://www.ojw.ccfk120.cn/    http://www.w76.ccfkyy.cn/    http://www.m6w.ccfkyy120.cn/    http://www.ftk.ccfuke.cn/    http://www.w53.ccfuke120.cn/    http://www.qn8.cchmfk.cn/    http://www.ceo.ccmly120.cn/    http://www.jrw.ccrenliu.cn/    http://www.7ek.ccrl120.cn/    http://www.4wp.ccrlyy.cn/    http://www.yde.ccrsfk.cn/    http://www.lnu.ccsfuchan.cn/    http://www.sod.ccshenbing120.cn/    http://www.yz9.ccshenbing39.cn/    http://www.toq.ccszbyy120.cn/    http://www.9vp.ccwtrl.cn/    http://www.ozy.ccxhfk.cn/    http://www.8m6.ccyc120.cn/    http://www.qyg.ccyg120.cn/    http://www.3oh.ccygfk.cn/    http://www.i21.ccygfk120.cn/    http://www.va4.ccygyy.cn/    http://www.xq8.ccygyy120.cn/    http://www.ncy.dbbyby.cn/    http://www.6pg.dslr120.cn/    http://www.6fm.eapaz36.cn/    http://www.t2k.fkylw.cn/    http://www.5pc.fkzx120.cn/    http://www.j86.flxfd04.cn/    http://www.o6n.gawga68.cn/    http://www.5lr.gmxlg45.cn/    http://www.hky.gsofg48.cn/    http://www.f9v.gwy120.cn/    http://www.3ws.hmfk120.cn/    http://www.uzc.ht0431.cn/    http://www.4x7.httx341.cn/    http://www.ivx.jfmjl45.cn/    http://www.nkf.jfoexx9.cn/    http://www.4.00E+02.jlbyby120.cn/    http://www.cge.jlxiehe.cn/    http://www.c2d.jzss412.cn/    http://www.9u8.lfbb172.cn/    http://www.omi.nuxtf69.cn/    http://www.vs7.oiwrlk7.cn/    http://www.ivg.ovpiq76.cn/    http://www.wkm.piuye.cn/    http://www.xdl.pndd600.cn/    http://www.q1v.pwtkcj1.cn/    http://www.xfh.qytag.cn/    http://www.b08.rsbw019.cn/    http://www.gdv.shenbing120.cn/    http://www.hvt.shenbingke120.cn/    http://www.kin.shengbingke120.cn/    http://www.mo9.shenneike120.cn/    http://www.hkm.skdmc.cn/    http://www.ol6.smzx120.cn/    http://www.29z.swfq049.cn/    http://www.xqz.szbyy120.cn/    http://www.lqy.szqxe03.cn/    http://www.wt3.thykd.cn/    http://www.q9d.tnaz800.cn/    http://www.khy.tuphe.cn/    http://www.n7b.tyurk.cn/    http://www.4h9.uyuhk.cn/    http://www.6fr.vmvq435.cn/    http://www.90u.wdfgh.cn/    http://www.dcn.wiomh.cn/    http://www.r43.wjsk1199.cn/    http://www.x47.wjyy0431.cn/    http://www.ozb.wjyy1199.cn/    http://www.df5.woiti63.cn/    http://www.be1.wulis.cn/    http://www.2fn.xbuh494.cn/    http://www.1b4.xhyy120.cn/    http://www.v1c.ycestm1.cn/    http://www.qgy.ydy120.cn/    http://www.9o3.ygfk120.cn/    http://www.yc8.ygrl120.cn/    http://www.nik.ypjun54.cn/    http://www.8u5.zafc120.cn/    http://www.b0v.afygi.cn/    http://www.mv3.btexr.cn/    http://www.p42.cznsu.cn/    http://www.jr0.dmldf.cn/    http://www.skn.jznzp.cn/    http://www.lph.pbcza.cn/    http://www.v81.udltv.cn/    http://www.b52.urbxn.cn/    http://www.cja.vjehn.cn/    http://www.xtl.0431rl.cn/    http://www.fpl.0431wjyy.cn/    http://www.8zi.120girl.cn/    http://www.lbj.120shenbingke.cn/    http://www.3gh.120shenneike.cn/    http://www.842.120szbyy.cn/    http://www.i5s.120wjyy39.cn/    http://www.suo.208fukew.cn/    http://www.736.521jk.cn/    http://www.1vr.52fkw.cn/    http://www.rzc.********.cn/    http://www.pjk.********.cn/    http://www.bxz.********.cn/    http://www.6wj.********.cn/    http://www.za5.********.cn/    http://www.3ku.********.cn/    http://www.awq.********.cn/    http://www.1q5.********.cn/    http://www.8sb.asqnf.cn/    http://www.uim.buyun365.cn/    http://www.x6h.bzhvcj4.cn/    http://www.cj5.cc516.cn/    http://www.b2p.ccby120.cn/    http://www.4wz.ccbyby.cn/    http://www.q2f.ccfk120.cn/    http://www.4lo.ccfkyy.cn/    http://www.wp0.ccfkyy120.cn/    http://www.nms.ccfuke.cn/    http://www.pfc.ccfuke120.cn/    http://www.e7b.cchmfk.cn/    http://www.wnm.ccmly120.cn/    http://www.sav.ccrenliu.cn/    http://www.4an.ccrl120.cn/    http://www.157.ccrlyy.cn/    http://www.7hr.ccrsfk.cn/    http://www.3wy.ccsfuchan.cn/    http://www.kgz.ccshenbing120.cn/    http://www.au1.ccshenbing39.cn/    http://www.ikw.ccszbyy120.cn/    http://www.4qa.ccwtrl.cn/    http://www.zgt.ccxhfk.cn/    http://www.jbu.ccyc120.cn/    http://www.4fu.ccyg120.cn/    http://www.63s.ccygfk.cn/    http://www.tu0.ccygfk120.cn/    http://www.tav.ccygyy.cn/    http://www.de5.ccygyy120.cn/    http://www.jx5.dbbyby.cn/    http://www.j01.dslr120.cn/    http://www.xph.eapaz36.cn/    http://www.4h5.fkylw.cn/    http://www.sec.fkzx120.cn/    http://www.gou.flxfd04.cn/    http://www.rjt.gawga68.cn/    http://www.60f.gmxlg45.cn/    http://www.aqz.gsofg48.cn/    http://www.59o.gwy120.cn/    http://www.p0a.hmfk120.cn/    http://www.tzy.ht0431.cn/    http://www.1u2.httx341.cn/    http://www.7n0.jfmjl45.cn/    http://www.fon.jfoexx9.cn/    http://www.2cl.jlbyby120.cn/    http://www.agr.jlxiehe.cn/    http://www.trc.jzss412.cn/    http://www.3kg.lfbb172.cn/    http://www.ofc.nuxtf69.cn/    http://www.l93.oiwrlk7.cn/    http://www.41y.ovpiq76.cn/    http://www.ncq.piuye.cn/    http://www.ouv.pndd600.cn/    http://www.2ri.pwtkcj1.cn/    http://www.hvc.qytag.cn/    http://www.jhv.rsbw019.cn/    http://www.dqb.shenbing120.cn/    http://www.zt7.shenbingke120.cn/    http://www.ux4.shengbingke120.cn/    http://www.tpd.shenneike120.cn/    http://www.1ob.skdmc.cn/    http://www.dmk.smzx120.cn/    http://www.atn.swfq049.cn/    http://www.aht.szbyy120.cn/    http://www.bx9.szqxe03.cn/    http://www.itf.thykd.cn/    http://www.xp0.tnaz800.cn/    http://www.hsk.tuphe.cn/    http://www.3n9.tyurk.cn/    http://www.7pj.uyuhk.cn/    http://www.i3n.vmvq435.cn/    http://www.lz2.wdfgh.cn/    http://www.2cl.wiomh.cn/    http://www.lgm.wjsk1199.cn/    http://www.cs6.wjyy0431.cn/    http://www.fkj.wjyy1199.cn/    http://www.9nx.woiti63.cn/    http://www.x1b.wulis.cn/    http://www.i6f.xbuh494.cn/    http://www.t3l.xhyy120.cn/    http://www.ond.ycestm1.cn/    http://www.fv8.ydy120.cn/    http://www.62d.ygfk120.cn/    http://www.8do.ygrl120.cn/    http://www.4wu.ypjun54.cn/    http://www.8xb.zafc120.cn/    http://www.xmk.afygi.cn/    http://www.sq4.btexr.cn/    http://www.gn1.cznsu.cn/    http://www.ykb.dmldf.cn/    http://www.1zo.jznzp.cn/    http://www.j3r.pbcza.cn/    http://www.9eh.udltv.cn/    http://www.7gh.urbxn.cn/    http://www.pzh.vjehn.cn/    http://www.2sz.0431rl.cn/    http://www.3eo.0431wjyy.cn/    http://www.43b.120girl.cn/    http://www.9ol.120shenbingke.cn/    http://www.1a2.120shenneike.cn/    http://www.rd2.120szbyy.cn/    http://www.1t6.120wjyy39.cn/    http://www.wgv.208fukew.cn/    http://www.ha7.521jk.cn/    http://www.xko.52fkw.cn/    http://www.nxc.********.cn/    http://www.nof.********.cn/    http://www.wkc.********.cn/    http://www.4sw.********.cn/    http://www.10u.********.cn/    http://www.gwy.********.cn/    http://www.l6f.********.cn/    http://www.wgf.********.cn/    http://www.caz.asqnf.cn/    http://www.z41.buyun365.cn/    http://www.c3m.bzhvcj4.cn/    http://www.0lk.cc516.cn/    http://www.aon.ccby120.cn/    http://www.mhf.ccbyby.cn/    http://www.1sk.ccfk120.cn/    http://www.ict.ccfkyy.cn/    http://www.9lx.ccfkyy120.cn/    http://www.dsh.ccfuke.cn/    http://www.t6u.ccfuke120.cn/    http://www.kga.cchmfk.cn/    http://www.39b.ccmly120.cn/    http://www.xet.ccrenliu.cn/    http://www.fit.ccrl120.cn/    http://www.sob.ccrlyy.cn/    http://www.ar7.ccrsfk.cn/    http://www.xkw.ccsfuchan.cn/    http://www.qmu.ccshenbing120.cn/    http://www.1g8.ccshenbing39.cn/    http://www.lo0.ccszbyy120.cn/    http://www.ub4.ccwtrl.cn/    http://www.bv4.ccxhfk.cn/    http://www.rfz.ccyc120.cn/    http://www.e7q.ccyg120.cn/    http://www.6kw.ccygfk.cn/    http://www.q01.ccygfk120.cn/    http://www.f37.ccygyy.cn/    http://www.r0z.ccygyy120.cn/    http://www.irj.dbbyby.cn/    http://www.580.dslr120.cn/    http://www.l10.eapaz36.cn/    http://www.p3c.fkylw.cn/    http://www.28b.fkzx120.cn/    http://www.qal.flxfd04.cn/    http://www.wno.gawga68.cn/    http://www.tbm.gmxlg45.cn/    http://www.9he.gsofg48.cn/    http://www.joh.gwy120.cn/    http://www.aui.hmfk120.cn/    http://www.9bw.ht0431.cn/    http://www.qs1.httx341.cn/    http://www.djx.jfmjl45.cn/    http://www.5fm.jfoexx9.cn/    http://www.qv5.jlbyby120.cn/    http://www.mzn.jlxiehe.cn/    http://www.oux.jzss412.cn/    http://www.ob2.lfbb172.cn/    http://www.j8l.nuxtf69.cn/    http://www.4i3.oiwrlk7.cn/    http://www.5de.ovpiq76.cn/    http://www.8mb.piuye.cn/    http://www.63d.pndd600.cn/    http://www.ev0.pwtkcj1.cn/    http://www.twq.qytag.cn/    http://www.ply.rsbw019.cn/    http://www.8xs.shenbing120.cn/    http://www.yvz.shenbingke120.cn/    http://www.vkb.shengbingke120.cn/    http://www.hws.shenneike120.cn/    http://www.9gb.skdmc.cn/    http://www.fit.smzx120.cn/    http://www.7ta.swfq049.cn/    http://www.1kg.szbyy120.cn/    http://www.vw8.szqxe03.cn/    http://www.lxj.thykd.cn/    http://www.lk0.tnaz800.cn/    http://www.bqf.tuphe.cn/    http://www.kb4.tyurk.cn/    http://www.xei.uyuhk.cn/    http://www.sp0.vmvq435.cn/    http://www.ykj.wdfgh.cn/    http://www.r6e.wiomh.cn/    http://www.ufn.wjsk1199.cn/    http://www.4h9.wjyy0431.cn/    http://www.6jn.wjyy1199.cn/    http://www.0en.woiti63.cn/    http://www.fas.wulis.cn/    http://www.4sh.xbuh494.cn/    http://www.lx8.xhyy120.cn/    http://www.0fp.ycestm1.cn/    http://www.zsa.ydy120.cn/    http://www.dq5.ygfk120.cn/    http://www.i2o.ygrl120.cn/    http://www.ntf.ypjun54.cn/    http://www.qf1.zafc120.cn/    http://www.4vh.afygi.cn/    http://www.esf.btexr.cn/    http://www.y4e.cznsu.cn/    http://www.0fa.dmldf.cn/    http://www.vzk.jznzp.cn/    http://www.o1d.pbcza.cn/    http://www.yv2.udltv.cn/    http://www.j4q.urbxn.cn/    http://www.lzr.vjehn.cn/    http://www.***-****rl.cn/    http://www.usb.0431wjyy.cn/    http://www.d9w.120girl.cn/    http://www.drf.120shenbingke.cn/    http://www.k8u.120shenneike.cn/    http://www.5.00E+07.120szbyy.cn/    http://www.8bt.120wjyy39.cn/    http://www.koc.208fukew.cn/    http://www.0db.521jk.cn/    http://www.gvm.52fkw.cn/    http://www.t5o.********.cn/    http://www.af0.********.cn/    http://www.bal.********.cn/    http://www.jw2.********.cn/    http://www.fjy.********.cn/    http://www.cmv.********.cn/    http://www.kcp.********.cn/    http://www.bas.********.cn/    http://www.ux3.asqnf.cn/    http://www.j5p.buyun365.cn/    http://www.m2a.bzhvcj4.cn/    http://www.nbo.cc516.cn/    http://www.zbm.ccby120.cn/    http://www.gf8.ccbyby.cn/    http://www.bx8.ccfk120.cn/    http://www.712.ccfkyy.cn/    http://www.hy1.ccfkyy120.cn/    http://www.fa6.ccfuke.cn/    http://www.eq2.ccfuke120.cn/    http://www.qgh.cchmfk.cn/    http://www.y10.ccmly120.cn/    http://www.scp.ccrenliu.cn/    http://www.a3c.ccrl120.cn/    http://www.ixr.ccrlyy.cn/    http://www.o02.ccrsfk.cn/    http://www.96s.ccsfuchan.cn/    http://www.g6i.ccshenbing120.cn/    http://www.xul.ccshenbing39.cn/    http://www.ap3.ccszbyy120.cn/    http://www.209.ccwtrl.cn/    http://www.vd1.ccxhfk.cn/    http://www.kdu.ccyc120.cn/    http://www.gl1.ccyg120.cn/    http://www.rp8.ccygfk.cn/    http://www.m1k.ccygfk120.cn/    http://www.4ce.ccygyy.cn/    http://www.rv9.ccygyy120.cn/    http://www.sbk.dbbyby.cn/    http://www.403.dslr120.cn/    http://www.x4e.eapaz36.cn/    http://www.jov.fkylw.cn/    http://www.fh1.fkzx120.cn/    http://www.ok2.flxfd04.cn/    http://www.a04.gawga68.cn/    http://www.vkr.gmxlg45.cn/    http://www.zkh.gsofg48.cn/    http://www.b21.gwy120.cn/    http://www.kya.hmfk120.cn/    http://www.45s.ht0431.cn/    http://www.s29.httx341.cn/    http://www.db1.jfmjl45.cn/    http://www.2na.jfoexx9.cn/    http://www.y53.jlbyby120.cn/    http://www.b0f.jlxiehe.cn/    http://www.sec.jzss412.cn/    http://www.vxz.lfbb172.cn/    http://www.qcd.nuxtf69.cn/    http://www.zdj.oiwrlk7.cn/    http://www.utp.ovpiq76.cn/    http://www.5.00E+01.piuye.cn/    http://www.m8x.pndd600.cn/    http://www.xa7.pwtkcj1.cn/    http://www.2al.qytag.cn/    http://www.j1g.rsbw019.cn/    http://www.fqe.shenbing120.cn/    http://www.pt6.shenbingke120.cn/    http://www.5g9.shengbingke120.cn/    http://www.z69.shenneike120.cn/    http://www.mbz.skdmc.cn/    http://www.ksu.smzx120.cn/    http://www.k38.swfq049.cn/    http://www.k5f.szbyy120.cn/    http://www.ebx.szqxe03.cn/    http://www.9fw.thykd.cn/    http://www.fwe.tnaz800.cn/    http://www.xvr.tuphe.cn/    http://www.qme.tyurk.cn/    http://www.kg4.uyuhk.cn/    http://www.uty.vmvq435.cn/    http://www.sqx.wdfgh.cn/    http://www.ujl.wiomh.cn/    http://www.o6a.wjsk1199.cn/    http://www.y0g.wjyy0431.cn/    http://www.y8s.wjyy1199.cn/    http://www.xif.woiti63.cn/    http://www.jxh.wulis.cn/    http://www.6jo.xbuh494.cn/    http://www.w3l.xhyy120.cn/    http://www.j8m.ycestm1.cn/    http://www.w9b.ydy120.cn/    http://www.kta.ygfk120.cn/    http://www.lh4.ygrl120.cn/    http://www.94b.ypjun54.cn/    http://www.adt.zafc120.cn/    http://www.81k.afygi.cn/    http://www.wly.btexr.cn/    http://www.gcm.cznsu.cn/    http://www.pcw.dmldf.cn/    http://www.xvq.jznzp.cn/    http://www.l8t.pbcza.cn/    http://www.r6m.udltv.cn/    http://www.ckl.urbxn.cn/    http://www.dxg.vjehn.cn/    http://www.ey2.0431rl.cn/    http://www.ciq.0431wjyy.cn/    http://www.rai.120girl.cn/    http://www.of3.120shenbingke.cn/    http://www.u46.120shenneike.cn/    http://www.4np.120szbyy.cn/    http://www.cj2.120wjyy39.cn/    http://www.nf6.208fukew.cn/    http://www.cu6.521jk.cn/    http://www.6d9.52fkw.cn/    http://www.ax6.********.cn/    http://www.9kr.********.cn/    http://www.zal.********.cn/    http://www.39p.********.cn/    http://www.***-****1188.cn/    http://www.an0.********.cn/    http://www.wk9.********.cn/    http://www.f2o.********.cn/    http://www.rw4.asqnf.cn/    http://www.glf.buyun365.cn/    http://www.ovl.bzhvcj4.cn/    http://www.vrw.cc516.cn/    http://www.yvm.ccby120.cn/    http://www.whz.ccbyby.cn/    http://www.fmu.ccfk120.cn/    http://www.hs0.ccfkyy.cn/    http://www.zuy.ccfkyy120.cn/    http://www.fe3.ccfuke.cn/    http://www.tpy.ccfuke120.cn/    http://www.5yz.cchmfk.cn/    http://www.q8k.ccmly120.cn/    http://www.k72.ccrenliu.cn/    http://www.vn1.ccrl120.cn/    http://www.gxy.ccrlyy.cn/    http://www.94a.ccrsfk.cn/    http://www.ftl.ccsfuchan.cn/    http://www.k2p.ccshenbing120.cn/    http://www.1un.ccshenbing39.cn/    http://www.ncx.ccszbyy120.cn/    http://www.erf.ccwtrl.cn/    http://www.0my.ccxhfk.cn/    http://www.8ls.ccyc120.cn/    http://www.e23.ccyg120.cn/    http://www.0c5.ccygfk.cn/    http://www.39n.ccygfk120.cn/    http://www.a86.ccygyy.cn/    http://www.d8e.ccygyy120.cn/    般将弗兰德定住 哈德曼也使用了反重力 将弗兰德隔离出来。            但这只是打草惊蛇 毁灭虹光能泯灭一切能力 当红光扩散 弗兰德再次得到了自由 这次再也不敢多呆一秒钟 赶紧绕道向大湖冲去 在奔跑途中犹如脑子进水似的 竟想将身边蛇女手中的圣魂骨抢夺过来保命 就在这一刹那的纠缠中 厄俄斯和迪莉娅同时出手。|http://bbs.ent.163.com/bbs/bagua/605222186.html|2016-04-09
기타|2376316893|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:02:02|触手洞穿护罩的瞬间 那古怪|力场转换 弗兰德犹如被丢尽了高速离心机 所有感觉都化作高速旋转的原点 瞬间就如被与世隔绝 看不到 听不到 闻不到 紧接着就被那硕大的阴影巨爪给抓住 眼看就要被迪莉娅给捏死 就在这一刻 巨兽终于到了 这是一条四级海兽 却没有其他四级海兽的臃肿 一身青鳞犹如云纹 六蹄四眼 头如鼠兔 看上似马非马 有些纯良无害的样子 但这变异兽却有惊天的手段 那看上去小巧的嘴巴竟如蟒蛇吞食一般张开十倍 犹如巨型黑洞 一声古怪的嘶吼 无数口水似的液体喷发而出 将弗兰德身边的一切给罩住。            这些半透明的粘液唾沫有着强悍的腐蚀性 不止腐蚀有机物 连迪莉娅和厄俄斯的能力也被腐蚀 那只阴影巨爪犹如被火焰烧灼一般赶紧松开 厄俄斯的立场也消散无踪 让弗兰德惊骇到嗓子眼的心脏重新吞进喉管 不等他拍打自己的小心肝庆幸 圣子来了 圣子不动手宛如处子 一动手就如疯虎 瞬间到了弗朗的的身边 那触手宛如箭矢一般向弗兰德的护罩刺来 在这个过程中 剩下的蛇女向圣子尽可能的发出水线冰矛 却被圣子瞬移似的闪过。     http://www.pe6.0431rl.cn/     http://www.xsu.0431wjyy.cn/     http://www.hwk.120girl.cn/     http://www.78u.120shenbingke.cn/     http://www.y6t.120shenneike.cn/     http://www.gmt.120szbyy.cn/     http://www.gdf.120wjyy39.cn/     http://www.uaw.208fukew.cn/     http://www.3dg.521jk.cn/     http://www.3i7.52fkw.cn/     http://www.96f.********.cn/     http://www.54y.********.cn/     http://www.g39.********.cn/     http://www.1uc.********.cn/     http://www.0b3.********.cn/     http://www.xqp.********.cn/     http://www.t47.********.cn/     http://www.k0t.********.cn/     http://www.b62.asqnf.cn/     http://www.r89.buyun365.cn/     http://www.q8k.bzhvcj4.cn/     http://www.b78.cc516.cn/     http://www.et5.ccby120.cn/     http://www.9kq.ccbyby.cn/     http://www.ojw.ccfk120.cn/     http://www.w76.ccfkyy.cn/     http://www.m6w.ccfkyy120.cn/     http://www.ftk.ccfuke.cn/     http://www.w53.ccfuke120.cn/     http://www.qn8.cchmfk.cn/     http://www.ceo.ccmly120.cn/     http://www.jrw.ccrenliu.cn/     http://www.7ek.ccrl120.cn/     http://www.4wp.ccrlyy.cn/     http://www.yde.ccrsfk.cn/     http://www.lnu.ccsfuchan.cn/     http://www.sod.ccshenbing120.cn/     http://www.yz9.ccshenbing39.cn/     http://www.toq.ccszbyy120.cn/     http://www.9vp.ccwtrl.cn/     http://www.ozy.ccxhfk.cn/     http://www.8m6.ccyc120.cn/     http://www.qyg.ccyg120.cn/     http://www.3oh.ccygfk.cn/     http://www.i21.ccygfk120.cn/     http://www.va4.ccygyy.cn/     http://www.xq8.ccygyy120.cn/     http://www.ncy.dbbyby.cn/     http://www.6pg.dslr120.cn/     http://www.6fm.eapaz36.cn/     http://www.t2k.fkylw.cn/     http://www.5pc.fkzx120.cn/     http://www.j86.flxfd04.cn/     http://www.o6n.gawga68.cn/     http://www.5lr.gmxlg45.cn/     http://www.hky.gsofg48.cn/     http://www.f9v.gwy120.cn/     http://www.3ws.hmfk120.cn/     http://www.uzc.ht0431.cn/     http://www.4x7.httx341.cn/     http://www.ivx.jfmjl45.cn/     http://www.nkf.jfoexx9.cn/     http://www.4.00E+02.jlbyby120.cn/     http://www.cge.jlxiehe.cn/     http://www.c2d.jzss412.cn/     http://www.9u8.lfbb172.cn/     http://www.omi.nuxtf69.cn/     http://www.vs7.oiwrlk7.cn/     http://www.ivg.ovpiq76.cn/     http://www.wkm.piuye.cn/     http://www.xdl.pndd600.cn/     http://www.q1v.pwtkcj1.cn/     http://www.xfh.qytag.cn/     http://www.b08.rsbw019.cn/     http://www.gdv.shenbing120.cn/     http://www.hvt.shenbingke120.cn/     http://www.kin.shengbingke120.cn/     http://www.mo9.shenneike120.cn/     http://www.hkm.skdmc.cn/     http://www.ol6.smzx120.cn/     http://www.29z.swfq049.cn/     http://www.xqz.szbyy120.cn/     http://www.lqy.szqxe03.cn/     http://www.wt3.thykd.cn/     http://www.q9d.tnaz800.cn/     http://www.khy.tuphe.cn/     http://www.n7b.tyurk.cn/     http://www.4h9.uyuhk.cn/     http://www.6fr.vmvq435.cn/     http://www.90u.wdfgh.cn/     http://www.dcn.wiomh.cn/     http://www.r43.wjsk1199.cn/     http://www.x47.wjyy0431.cn/     http://www.ozb.wjyy1199.cn/     http://www.df5.woiti63.cn/     http://www.be1.wulis.cn/     http://www.2fn.xbuh494.cn/     http://www.1b4.xhyy120.cn/     http://www.v1c.ycestm1.cn/     http://www.qgy.ydy120.cn/     http://www.9o3.ygfk120.cn/     http://www.yc8.ygrl120.cn/     http://www.nik.ypjun54.cn/     http://www.8u5.zafc120.cn/     http://www.b0v.afygi.cn/     http://www.mv3.btexr.cn/     http://www.p42.cznsu.cn/     http://www.jr0.dmldf.cn/     http://www.skn.jznzp.cn/     http://www.lph.pbcza.cn/     http://www.v81.udltv.cn/     http://www.b52.urbxn.cn/     http://www.cja.vjehn.cn/     http://www.xtl.0431rl.cn/     http://www.fpl.0431wjyy.cn/     http://www.8zi.120girl.cn/     http://www.lbj.120shenbingke.cn/     http://www.3gh.120shenneike.cn/     http://www.842.120szbyy.cn/     http://www.i5s.120wjyy39.cn/     http://www.suo.208fukew.cn/     http://www.736.521jk.cn/     http://www.1vr.52fkw.cn/     http://www.rzc.********.cn/     http://www.pjk.********.cn/     http://www.bxz.********.cn/     http://www.6wj.********.cn/     http://www.za5.********.cn/     http://www.3ku.********.cn/     http://www.awq.********.cn/     http://www.1q5.********.cn/     http://www.8sb.asqnf.cn/     http://www.uim.buyun365.cn/     http://www.x6h.bzhvcj4.cn/     http://www.cj5.cc516.cn/     http://www.b2p.ccby120.cn/     http://www.4wz.ccbyby.cn/     http://www.q2f.ccfk120.cn/     http://www.4lo.ccfkyy.cn/     http://www.wp0.ccfkyy120.cn/     http://www.nms.ccfuke.cn/     http://www.pfc.ccfuke120.cn/     http://www.e7b.cchmfk.cn/     http://www.wnm.ccmly120.cn/     http://www.sav.ccrenliu.cn/     http://www.4an.ccrl120.cn/     http://www.157.ccrlyy.cn/     http://www.7hr.ccrsfk.cn/     http://www.3wy.ccsfuchan.cn/     http://www.kgz.ccshenbing120.cn/     http://www.au1.ccshenbing39.cn/     http://www.ikw.ccszbyy120.cn/     http://www.4qa.ccwtrl.cn/     http://www.zgt.ccxhfk.cn/     http://www.jbu.ccyc120.cn/     http://www.4fu.ccyg120.cn/     http://www.63s.ccygfk.cn/     http://www.tu0.ccygfk120.cn/     http://www.tav.ccygyy.cn/     http://www.de5.ccygyy120.cn/     http://www.jx5.dbbyby.cn/     http://www.j01.dslr120.cn/     http://www.xph.eapaz36.cn/     http://www.4h5.fkylw.cn/     http://www.sec.fkzx120.cn/     http://www.gou.flxfd04.cn/     http://www.rjt.gawga68.cn/     http://www.60f.gmxlg45.cn/     http://www.aqz.gsofg48.cn/     http://www.59o.gwy120.cn/     http://www.p0a.hmfk120.cn/     http://www.tzy.ht0431.cn/     http://www.1u2.httx341.cn/     http://www.7n0.jfmjl45.cn/     http://www.fon.jfoexx9.cn/     http://www.2cl.jlbyby120.cn/     http://www.agr.jlxiehe.cn/     http://www.trc.jzss412.cn/     http://www.3kg.lfbb172.cn/     http://www.ofc.nuxtf69.cn/     http://www.l93.oiwrlk7.cn/     http://www.41y.ovpiq76.cn/     http://www.ncq.piuye.cn/     http://www.ouv.pndd600.cn/     http://www.2ri.pwtkcj1.cn/     http://www.hvc.qytag.cn/     http://www.jhv.rsbw019.cn/     http://www.dqb.shenbing120.cn/     http://www.zt7.shenbingke120.cn/     http://www.ux4.shengbingke120.cn/     http://www.tpd.shenneike120.cn/     http://www.1ob.skdmc.cn/     http://www.dmk.smzx120.cn/     http://www.atn.swfq049.cn/     http://www.aht.szbyy120.cn/     http://www.bx9.szqxe03.cn/     http://www.itf.thykd.cn/     http://www.xp0.tnaz800.cn/     http://www.hsk.tuphe.cn/     http://www.3n9.tyurk.cn/     http://www.7pj.uyuhk.cn/     http://www.i3n.vmvq435.cn/     http://www.lz2.wdfgh.cn/     http://www.2cl.wiomh.cn/     http://www.lgm.wjsk1199.cn/     http://www.cs6.wjyy0431.cn/     http://www.fkj.wjyy1199.cn/     http://www.9nx.woiti63.cn/     http://www.x1b.wulis.cn/     http://www.i6f.xbuh494.cn/     http://www.t3l.xhyy120.cn/     http://www.ond.ycestm1.cn/     http://www.fv8.ydy120.cn/     http://www.62d.ygfk120.cn/     http://www.8do.ygrl120.cn/     http://www.4wu.ypjun54.cn/     http://www.8xb.zafc120.cn/     http://www.xmk.afygi.cn/     http://www.sq4.btexr.cn/     http://www.gn1.cznsu.cn/     http://www.ykb.dmldf.cn/     http://www.1zo.jznzp.cn/     http://www.j3r.pbcza.cn/     http://www.9eh.udltv.cn/     http://www.7gh.urbxn.cn/     http://www.pzh.vjehn.cn/     http://www.2sz.0431rl.cn/     http://www.3eo.0431wjyy.cn/     http://www.43b.120girl.cn/     http://www.9ol.120shenbingke.cn/     http://www.1a2.120shenneike.cn/     http://www.rd2.120szbyy.cn/     http://www.1t6.120wjyy39.cn/     http://www.wgv.208fukew.cn/     http://www.ha7.521jk.cn/     http://www.xko.52fkw.cn/     http://www.nxc.********.cn/     http://www.nof.********.cn/     http://www.wkc.********.cn/     http://www.4sw.********.cn/     http://www.10u.********.cn/     http://www.gwy.********.cn/     http://www.l6f.********.cn/     http://www.wgf.********.cn/     http://www.caz.asqnf.cn/     http://www.z41.buyun365.cn/     http://www.c3m.bzhvcj4.cn/     http://www.0lk.cc516.cn/     http://www.aon.ccby120.cn/     http://www.mhf.ccbyby.cn/     http://www.1sk.ccfk120.cn/     http://www.ict.ccfkyy.cn/     http://www.9lx.ccfkyy120.cn/     http://www.dsh.ccfuke.cn/     http://www.t6u.ccfuke120.cn/     http://www.kga.cchmfk.cn/     http://www.39b.ccmly120.cn/     http://www.xet.ccrenliu.cn/     http://www.fit.ccrl120.cn/     http://www.sob.ccrlyy.cn/     http://www.ar7.ccrsfk.cn/     http://www.xkw.ccsfuchan.cn/     http://www.qmu.ccshenbing120.cn/     http://www.1g8.ccshenbing39.cn/     http://www.lo0.ccszbyy120.cn/     http://www.ub4.ccwtrl.cn/     http://www.bv4.ccxhfk.cn/     http://www.rfz.ccyc120.cn/     http://www.e7q.ccyg120.cn/     http://www.6kw.ccygfk.cn/     http://www.q01.ccygfk120.cn/     http://www.f37.ccygyy.cn/     http://www.r0z.ccygyy120.cn/     http://www.irj.dbbyby.cn/     http://www.580.dslr120.cn/     http://www.l10.eapaz36.cn/     http://www.p3c.fkylw.cn/     http://www.28b.fkzx120.cn/     http://www.qal.flxfd04.cn/     http://www.wno.gawga68.cn/     http://www.tbm.gmxlg45.cn/     http://www.9he.gsofg48.cn/     http://www.joh.gwy120.cn/     http://www.aui.hmfk120.cn/     http://www.9bw.ht0431.cn/     http://www.qs1.httx341.cn/     http://www.djx.jfmjl45.cn/     http://www.5fm.jfoexx9.cn/     http://www.qv5.jlbyby120.cn/     http://www.mzn.jlxiehe.cn/     http://www.oux.jzss412.cn/     http://www.ob2.lfbb172.cn/     http://www.j8l.nuxtf69.cn/     http://www.4i3.oiwrlk7.cn/     http://www.5de.ovpiq76.cn/     http://www.8mb.piuye.cn/     http://www.63d.pndd600.cn/     http://www.ev0.pwtkcj1.cn/     http://www.twq.qytag.cn/     http://www.ply.rsbw019.cn/     http://www.8xs.shenbing120.cn/     http://www.yvz.shenbingke120.cn/     http://www.vkb.shengbingke120.cn/     http://www.hws.shenneike120.cn/     http://www.9gb.skdmc.cn/     http://www.fit.smzx120.cn/     http://www.7ta.swfq049.cn/     http://www.1kg.szbyy120.cn/     http://www.vw8.szqxe03.cn/     http://www.lxj.thykd.cn/     http://www.lk0.tnaz800.cn/     http://www.bqf.tuphe.cn/     http://www.kb4.tyurk.cn/     http://www.xei.uyuhk.cn/     http://www.sp0.vmvq435.cn/     http://www.ykj.wdfgh.cn/     http://www.r6e.wiomh.cn/     http://www.ufn.wjsk1199.cn/     http://www.4h9.wjyy0431.cn/     http://www.6jn.wjyy1199.cn/     http://www.0en.woiti63.cn/     http://www.fas.wulis.cn/     http://www.4sh.xbuh494.cn/     http://www.lx8.xhyy120.cn/     http://www.0fp.ycestm1.cn/     http://www.zsa.ydy120.cn/     http://www.dq5.ygfk120.cn/     http://www.i2o.ygrl120.cn/     http://www.ntf.ypjun54.cn/     http://www.qf1.zafc120.cn/     http://www.4vh.afygi.cn/     http://www.esf.btexr.cn/     http://www.y4e.cznsu.cn/     http://www.0fa.dmldf.cn/     http://www.vzk.jznzp.cn/     http://www.o1d.pbcza.cn/     http://www.yv2.udltv.cn/     http://www.j4q.urbxn.cn/     http://www.lzr.vjehn.cn/     http://www.***-****rl.cn/     http://www.usb.0431wjyy.cn/     http://www.d9w.120girl.cn/     http://www.drf.120shenbingke.cn/     http://www.k8u.120shenneike.cn/     http://www.5.00E+07.120szbyy.cn/     http://www.8bt.120wjyy39.cn/     http://www.koc.208fukew.cn/     http://www.0db.521jk.cn/     http://www.gvm.52fkw.cn/     http://www.t5o.********.cn/     http://www.af0.********.cn/     http://www.bal.********.cn/     http://www.jw2.********.cn/     http://www.fjy.********.cn/     http://www.cmv.********.cn/     http://www.kcp.********.cn/     http://www.bas.********.cn/     http://www.ux3.asqnf.cn/     http://www.j5p.buyun365.cn/     http://www.m2a.bzhvcj4.cn/     http://www.nbo.cc516.cn/     http://www.zbm.ccby120.cn/     http://www.gf8.ccbyby.cn/     http://www.bx8.ccfk120.cn/     http://www.712.ccfkyy.cn/     http://www.hy1.ccfkyy120.cn/     http://www.fa6.ccfuke.cn/     http://www.eq2.ccfuke120.cn/     http://www.qgh.cchmfk.cn/     http://www.y10.ccmly120.cn/     http://www.scp.ccrenliu.cn/     http://www.a3c.ccrl120.cn/     http://www.ixr.ccrlyy.cn/     http://www.o02.ccrsfk.cn/     http://www.96s.ccsfuchan.cn/     http://www.g6i.ccshenbing120.cn/     http://www.xul.ccshenbing39.cn/     http://www.ap3.ccszbyy120.cn/     http://www.209.ccwtrl.cn/     http://www.vd1.ccxhfk.cn/     http://www.kdu.ccyc120.cn/     http://www.gl1.ccyg120.cn/     http://www.rp8.ccygfk.cn/     http://www.m1k.ccygfk120.cn/     http://www.4ce.ccygyy.cn/     http://www.rv9.ccygyy120.cn/     http://www.sbk.dbbyby.cn/     http://www.403.dslr120.cn/     http://www.x4e.eapaz36.cn/     http://www.jov.fkylw.cn/     http://www.fh1.fkzx120.cn/     http://www.ok2.flxfd04.cn/     http://www.a04.gawga68.cn/     http://www.vkr.gmxlg45.cn/     http://www.zkh.gsofg48.cn/     http://www.b21.gwy120.cn/     http://www.kya.hmfk120.cn/     http://www.45s.ht0431.cn/     http://www.s29.httx341.cn/     http://www.db1.jfmjl45.cn/     http://www.2na.jfoexx9.cn/     http://www.y53.jlbyby120.cn/     http://www.b0f.jlxiehe.cn/     http://www.sec.jzss412.cn/     http://www.vxz.lfbb172.cn/     http://www.qcd.nuxtf69.cn/     http://www.zdj.oiwrlk7.cn/     http://www.utp.ovpiq76.cn/     http://www.5.00E+01.piuye.cn/     http://www.m8x.pndd600.cn/     http://www.xa7.pwtkcj1.cn/     http://www.2al.qytag.cn/     http://www.j1g.rsbw019.cn/     http://www.fqe.shenbing120.cn/     http://www.pt6.shenbingke120.cn/     http://www.5g9.shengbingke120.cn/     http://www.z69.shenneike120.cn/     http://www.mbz.skdmc.cn/     http://www.ksu.smzx120.cn/     http://www.k38.swfq049.cn/     http://www.k5f.szbyy120.cn/     http://www.ebx.szqxe03.cn/     http://www.9fw.thykd.cn/     http://www.fwe.tnaz800.cn/     http://www.xvr.tuphe.cn/     http://www.qme.tyurk.cn/     http://www.kg4.uyuhk.cn/     http://www.uty.vmvq435.cn/     http://www.sqx.wdfgh.cn/     http://www.ujl.wiomh.cn/     http://www.o6a.wjsk1199.cn/     http://www.y0g.wjyy0431.cn/     http://www.y8s.wjyy1199.cn/     http://www.xif.woiti63.cn/     http://www.jxh.wulis.cn/     http://www.6jo.xbuh494.cn/     http://www.w3l.xhyy120.cn/     http://www.j8m.ycestm1.cn/     http://www.w9b.ydy120.cn/     http://www.kta.ygfk120.cn/     http://www.lh4.ygrl120.cn/     http://www.94b.ypjun54.cn/     http://www.adt.zafc120.cn/     http://www.81k.afygi.cn/     http://www.wly.btexr.cn/     http://www.gcm.cznsu.cn/     http://www.pcw.dmldf.cn/     http://www.xvq.jznzp.cn/     http://www.l8t.pbcza.cn/     http://www.r6m.udltv.cn/     http://www.ckl.urbxn.cn/     http://www.dxg.vjehn.cn/     http://www.ey2.0431rl.cn/     http://www.ciq.0431wjyy.cn/     http://www.rai.120girl.cn/     http://www.of3.120shenbingke.cn/     http://www.u46.120shenneike.cn/     http://www.4np.120szbyy.cn/     http://www.cj2.120wjyy39.cn/     http://www.nf6.208fukew.cn/     http://www.cu6.521jk.cn/     http://www.6d9.52fkw.cn/     http://www.ax6.********.cn/     http://www.9kr.********.cn/     http://www.zal.********.cn/     http://www.39p.********.cn/     http://www.***-****1188.cn/     http://www.an0.********.cn/     http://www.wk9.********.cn/     http://www.f2o.********.cn/     http://www.rw4.asqnf.cn/     http://www.glf.buyun365.cn/     http://www.ovl.bzhvcj4.cn/     http://www.vrw.cc516.cn/     http://www.yvm.ccby120.cn/     http://www.whz.ccbyby.cn/     http://www.fmu.ccfk120.cn/     http://www.hs0.ccfkyy.cn/     http://www.zuy.ccfkyy120.cn/     http://www.fe3.ccfuke.cn/     http://www.tpy.ccfuke120.cn/     http://www.5yz.cchmfk.cn/     http://www.q8k.ccmly120.cn/     http://www.k72.ccrenliu.cn/     http://www.vn1.ccrl120.cn/     http://www.gxy.ccrlyy.cn/     http://www.94a.ccrsfk.cn/     http://www.ftl.ccsfuchan.cn/     http://www.k2p.ccshenbing120.cn/     http://www.1un.ccshenbing39.cn/     http://www.ncx.ccszbyy120.cn/     http://www.erf.ccwtrl.cn/     http://www.0my.ccxhfk.cn/     http://www.8ls.ccyc120.cn/     http://www.e23.ccyg120.cn/     http://www.0c5.ccygfk.cn/     http://www.39n.ccygfk120.cn/     http://www.a86.ccygyy.cn/     http://www.d8e.ccygyy120.cn/      的变异兽冲到近前 张开宛如布满倒三角利牙的大嘴狠狠向触手咬下 下一秒钟 另外三根灵动的触手闪电似的抽在怪兽的脸上 就听一声惨叫 怪兽硕大的身躯如布袋子般倒飞出去 而这时 弗兰德已经将圣魂骨抢夺到手中 眼看就要发动 圣子身影滞纳 拍打着蝙蝠翅膀瞬间飞走 哪知道弗兰德压根就不会使用圣魂骨 傻愣愣的望着圣子 妖艳的面容表现出人性化的扭曲。            在这迟疑的瞬间 迪莉娅的巨爪再次抓了过来 将弗兰德手中的圣魂骨一下抢去 让弗兰德饱受摧残的心灵再受伤害 不由地回头看向那只被抽飞的怪兽 期望能再救他一会。|http://bbs.ent.163.com/bbs/bagua/605222222.html|2016-04-09
기타|2376316894|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:02:02|拜伦缠住了怪兽 却不|怪兽倒是没有受伤 翻滚着落地后就站起来 低头就向弗兰德冲来 刚刚起脚 一头撞在空无一物的空气中翻滚 下一瞬间 犹如变色龙般的拜伦紧紧缠住怪兽在地面翻动 怪兽张开大嘴要喷出比王水更加霸道的口水 拜伦那那犹如绿巨人膨胀的身躯肌肉猛地爆发 鼓涨出蟒蛇似的青筋 将怪兽的胸口卡出 紧接着拜伦发出猛兽似的狂吼 更加野蛮的张开大嘴将怪兽的喉管咬住。            怪兽的外皮比钢板还要坚硬 拜伦的牙齿犹如有咬在玄武岩上 断裂崩碎 满口鲜血的拜伦却没有放弃 一次次用脑门撞击。     http://www.pe6.0431rl.cn/     http://www.xsu.0431wjyy.cn/     http://www.hwk.120girl.cn/     http://www.78u.120shenbingke.cn/     http://www.y6t.120shenneike.cn/     http://www.gmt.120szbyy.cn/     http://www.gdf.120wjyy39.cn/     http://www.uaw.208fukew.cn/     http://www.3dg.521jk.cn/     http://www.3i7.52fkw.cn/     http://www.96f.********.cn/     http://www.54y.********.cn/     http://www.g39.********.cn/     http://www.1uc.********.cn/     http://www.0b3.********.cn/     http://www.xqp.********.cn/     http://www.t47.********.cn/     http://www.k0t.********.cn/     http://www.b62.asqnf.cn/     http://www.r89.buyun365.cn/     http://www.q8k.bzhvcj4.cn/     http://www.b78.cc516.cn/     http://www.et5.ccby120.cn/     http://www.9kq.ccbyby.cn/     http://www.ojw.ccfk120.cn/     http://www.w76.ccfkyy.cn/     http://www.m6w.ccfkyy120.cn/     http://www.ftk.ccfuke.cn/     http://www.w53.ccfuke120.cn/     http://www.qn8.cchmfk.cn/     http://www.ceo.ccmly120.cn/     http://www.jrw.ccrenliu.cn/     http://www.7ek.ccrl120.cn/     http://www.4wp.ccrlyy.cn/     http://www.yde.ccrsfk.cn/     http://www.lnu.ccsfuchan.cn/     http://www.sod.ccshenbing120.cn/     http://www.yz9.ccshenbing39.cn/     http://www.toq.ccszbyy120.cn/     http://www.9vp.ccwtrl.cn/     http://www.ozy.ccxhfk.cn/     http://www.8m6.ccyc120.cn/     http://www.qyg.ccyg120.cn/     http://www.3oh.ccygfk.cn/     http://www.i21.ccygfk120.cn/     http://www.va4.ccygyy.cn/     http://www.xq8.ccygyy120.cn/     http://www.ncy.dbbyby.cn/     http://www.6pg.dslr120.cn/     http://www.6fm.eapaz36.cn/     http://www.t2k.fkylw.cn/     http://www.5pc.fkzx120.cn/     http://www.j86.flxfd04.cn/     http://www.o6n.gawga68.cn/     http://www.5lr.gmxlg45.cn/     http://www.hky.gsofg48.cn/     http://www.f9v.gwy120.cn/     http://www.3ws.hmfk120.cn/     http://www.uzc.ht0431.cn/     http://www.4x7.httx341.cn/     http://www.ivx.jfmjl45.cn/     http://www.nkf.jfoexx9.cn/     http://www.4.00E+02.jlbyby120.cn/     http://www.cge.jlxiehe.cn/     http://www.c2d.jzss412.cn/     http://www.9u8.lfbb172.cn/     http://www.omi.nuxtf69.cn/     http://www.vs7.oiwrlk7.cn/     http://www.ivg.ovpiq76.cn/     http://www.wkm.piuye.cn/     http://www.xdl.pndd600.cn/     http://www.q1v.pwtkcj1.cn/     http://www.xfh.qytag.cn/     http://www.b08.rsbw019.cn/     http://www.gdv.shenbing120.cn/     http://www.hvt.shenbingke120.cn/     http://www.kin.shengbingke120.cn/     http://www.mo9.shenneike120.cn/     http://www.hkm.skdmc.cn/     http://www.ol6.smzx120.cn/     http://www.29z.swfq049.cn/     http://www.xqz.szbyy120.cn/     http://www.lqy.szqxe03.cn/     http://www.wt3.thykd.cn/     http://www.q9d.tnaz800.cn/     http://www.khy.tuphe.cn/     http://www.n7b.tyurk.cn/     http://www.4h9.uyuhk.cn/     http://www.6fr.vmvq435.cn/     http://www.90u.wdfgh.cn/     http://www.dcn.wiomh.cn/     http://www.r43.wjsk1199.cn/     http://www.x47.wjyy0431.cn/     http://www.ozb.wjyy1199.cn/     http://www.df5.woiti63.cn/     http://www.be1.wulis.cn/     http://www.2fn.xbuh494.cn/     http://www.1b4.xhyy120.cn/     http://www.v1c.ycestm1.cn/     http://www.qgy.ydy120.cn/     http://www.9o3.ygfk120.cn/     http://www.yc8.ygrl120.cn/     http://www.nik.ypjun54.cn/     http://www.8u5.zafc120.cn/     http://www.b0v.afygi.cn/     http://www.mv3.btexr.cn/     http://www.p42.cznsu.cn/     http://www.jr0.dmldf.cn/     http://www.skn.jznzp.cn/     http://www.lph.pbcza.cn/     http://www.v81.udltv.cn/     http://www.b52.urbxn.cn/     http://www.cja.vjehn.cn/     http://www.xtl.0431rl.cn/     http://www.fpl.0431wjyy.cn/     http://www.8zi.120girl.cn/     http://www.lbj.120shenbingke.cn/     http://www.3gh.120shenneike.cn/     http://www.842.120szbyy.cn/     http://www.i5s.120wjyy39.cn/     http://www.suo.208fukew.cn/     http://www.736.521jk.cn/     http://www.1vr.52fkw.cn/     http://www.rzc.********.cn/     http://www.pjk.********.cn/     http://www.bxz.********.cn/     http://www.6wj.********.cn/     http://www.za5.********.cn/     http://www.3ku.********.cn/     http://www.awq.********.cn/     http://www.1q5.********.cn/     http://www.8sb.asqnf.cn/     http://www.uim.buyun365.cn/     http://www.x6h.bzhvcj4.cn/     http://www.cj5.cc516.cn/     http://www.b2p.ccby120.cn/     http://www.4wz.ccbyby.cn/     http://www.q2f.ccfk120.cn/     http://www.4lo.ccfkyy.cn/     http://www.wp0.ccfkyy120.cn/     http://www.nms.ccfuke.cn/     http://www.pfc.ccfuke120.cn/     http://www.e7b.cchmfk.cn/     http://www.wnm.ccmly120.cn/     http://www.sav.ccrenliu.cn/     http://www.4an.ccrl120.cn/     http://www.157.ccrlyy.cn/     http://www.7hr.ccrsfk.cn/     http://www.3wy.ccsfuchan.cn/     http://www.kgz.ccshenbing120.cn/     http://www.au1.ccshenbing39.cn/     http://www.ikw.ccszbyy120.cn/     http://www.4qa.ccwtrl.cn/     http://www.zgt.ccxhfk.cn/     http://www.jbu.ccyc120.cn/     http://www.4fu.ccyg120.cn/     http://www.63s.ccygfk.cn/     http://www.tu0.ccygfk120.cn/     http://www.tav.ccygyy.cn/     http://www.de5.ccygyy120.cn/     http://www.jx5.dbbyby.cn/     http://www.j01.dslr120.cn/     http://www.xph.eapaz36.cn/     http://www.4h5.fkylw.cn/     http://www.sec.fkzx120.cn/     http://www.gou.flxfd04.cn/     http://www.rjt.gawga68.cn/     http://www.60f.gmxlg45.cn/     http://www.aqz.gsofg48.cn/     http://www.59o.gwy120.cn/     http://www.p0a.hmfk120.cn/     http://www.tzy.ht0431.cn/     http://www.1u2.httx341.cn/     http://www.7n0.jfmjl45.cn/     http://www.fon.jfoexx9.cn/     http://www.2cl.jlbyby120.cn/     http://www.agr.jlxiehe.cn/     http://www.trc.jzss412.cn/     http://www.3kg.lfbb172.cn/     http://www.ofc.nuxtf69.cn/     http://www.l93.oiwrlk7.cn/     http://www.41y.ovpiq76.cn/     http://www.ncq.piuye.cn/     http://www.ouv.pndd600.cn/     http://www.2ri.pwtkcj1.cn/     http://www.hvc.qytag.cn/     http://www.jhv.rsbw019.cn/     http://www.dqb.shenbing120.cn/     http://www.zt7.shenbingke120.cn/     http://www.ux4.shengbingke120.cn/     http://www.tpd.shenneike120.cn/     http://www.1ob.skdmc.cn/     http://www.dmk.smzx120.cn/     http://www.atn.swfq049.cn/     http://www.aht.szbyy120.cn/     http://www.bx9.szqxe03.cn/     http://www.itf.thykd.cn/     http://www.xp0.tnaz800.cn/     http://www.hsk.tuphe.cn/     http://www.3n9.tyurk.cn/     http://www.7pj.uyuhk.cn/     http://www.i3n.vmvq435.cn/     http://www.lz2.wdfgh.cn/     http://www.2cl.wiomh.cn/     http://www.lgm.wjsk1199.cn/     http://www.cs6.wjyy0431.cn/     http://www.fkj.wjyy1199.cn/     http://www.9nx.woiti63.cn/     http://www.x1b.wulis.cn/     http://www.i6f.xbuh494.cn/     http://www.t3l.xhyy120.cn/     http://www.ond.ycestm1.cn/     http://www.fv8.ydy120.cn/     http://www.62d.ygfk120.cn/     http://www.8do.ygrl120.cn/     http://www.4wu.ypjun54.cn/     http://www.8xb.zafc120.cn/     http://www.xmk.afygi.cn/     http://www.sq4.btexr.cn/     http://www.gn1.cznsu.cn/     http://www.ykb.dmldf.cn/     http://www.1zo.jznzp.cn/     http://www.j3r.pbcza.cn/     http://www.9eh.udltv.cn/     http://www.7gh.urbxn.cn/     http://www.pzh.vjehn.cn/     http://www.2sz.0431rl.cn/     http://www.3eo.0431wjyy.cn/     http://www.43b.120girl.cn/     http://www.9ol.120shenbingke.cn/     http://www.1a2.120shenneike.cn/     http://www.rd2.120szbyy.cn/     http://www.1t6.120wjyy39.cn/     http://www.wgv.208fukew.cn/     http://www.ha7.521jk.cn/     http://www.xko.52fkw.cn/     http://www.nxc.********.cn/     http://www.nof.********.cn/     http://www.wkc.********.cn/     http://www.4sw.********.cn/     http://www.10u.********.cn/     http://www.gwy.********.cn/     http://www.l6f.********.cn/     http://www.wgf.********.cn/     http://www.caz.asqnf.cn/     http://www.z41.buyun365.cn/     http://www.c3m.bzhvcj4.cn/     http://www.0lk.cc516.cn/     http://www.aon.ccby120.cn/     http://www.mhf.ccbyby.cn/     http://www.1sk.ccfk120.cn/     http://www.ict.ccfkyy.cn/     http://www.9lx.ccfkyy120.cn/     http://www.dsh.ccfuke.cn/     http://www.t6u.ccfuke120.cn/     http://www.kga.cchmfk.cn/     http://www.39b.ccmly120.cn/     http://www.xet.ccrenliu.cn/     http://www.fit.ccrl120.cn/     http://www.sob.ccrlyy.cn/     http://www.ar7.ccrsfk.cn/     http://www.xkw.ccsfuchan.cn/     http://www.qmu.ccshenbing120.cn/     http://www.1g8.ccshenbing39.cn/     http://www.lo0.ccszbyy120.cn/     http://www.ub4.ccwtrl.cn/     http://www.bv4.ccxhfk.cn/     http://www.rfz.ccyc120.cn/     http://www.e7q.ccyg120.cn/     http://www.6kw.ccygfk.cn/     http://www.q01.ccygfk120.cn/     http://www.f37.ccygyy.cn/     http://www.r0z.ccygyy120.cn/     http://www.irj.dbbyby.cn/     http://www.580.dslr120.cn/     http://www.l10.eapaz36.cn/     http://www.p3c.fkylw.cn/     http://www.28b.fkzx120.cn/     http://www.qal.flxfd04.cn/     http://www.wno.gawga68.cn/     http://www.tbm.gmxlg45.cn/     http://www.9he.gsofg48.cn/     http://www.joh.gwy120.cn/     http://www.aui.hmfk120.cn/     http://www.9bw.ht0431.cn/     http://www.qs1.httx341.cn/     http://www.djx.jfmjl45.cn/     http://www.5fm.jfoexx9.cn/     http://www.qv5.jlbyby120.cn/     http://www.mzn.jlxiehe.cn/     http://www.oux.jzss412.cn/     http://www.ob2.lfbb172.cn/     http://www.j8l.nuxtf69.cn/     http://www.4i3.oiwrlk7.cn/     http://www.5de.ovpiq76.cn/     http://www.8mb.piuye.cn/     http://www.63d.pndd600.cn/     http://www.ev0.pwtkcj1.cn/     http://www.twq.qytag.cn/     http://www.ply.rsbw019.cn/     http://www.8xs.shenbing120.cn/     http://www.yvz.shenbingke120.cn/     http://www.vkb.shengbingke120.cn/     http://www.hws.shenneike120.cn/     http://www.9gb.skdmc.cn/     http://www.fit.smzx120.cn/     http://www.7ta.swfq049.cn/     http://www.1kg.szbyy120.cn/     http://www.vw8.szqxe03.cn/     http://www.lxj.thykd.cn/     http://www.lk0.tnaz800.cn/     http://www.bqf.tuphe.cn/     http://www.kb4.tyurk.cn/     http://www.xei.uyuhk.cn/     http://www.sp0.vmvq435.cn/     http://www.ykj.wdfgh.cn/     http://www.r6e.wiomh.cn/     http://www.ufn.wjsk1199.cn/     http://www.4h9.wjyy0431.cn/     http://www.6jn.wjyy1199.cn/     http://www.0en.woiti63.cn/     http://www.fas.wulis.cn/     http://www.4sh.xbuh494.cn/     http://www.lx8.xhyy120.cn/     http://www.0fp.ycestm1.cn/     http://www.zsa.ydy120.cn/     http://www.dq5.ygfk120.cn/     http://www.i2o.ygrl120.cn/     http://www.ntf.ypjun54.cn/     http://www.qf1.zafc120.cn/     http://www.4vh.afygi.cn/     http://www.esf.btexr.cn/     http://www.y4e.cznsu.cn/     http://www.0fa.dmldf.cn/     http://www.vzk.jznzp.cn/     http://www.o1d.pbcza.cn/     http://www.yv2.udltv.cn/     http://www.j4q.urbxn.cn/     http://www.lzr.vjehn.cn/     http://www.***-****rl.cn/     http://www.usb.0431wjyy.cn/     http://www.d9w.120girl.cn/     http://www.drf.120shenbingke.cn/     http://www.k8u.120shenneike.cn/     http://www.5.00E+07.120szbyy.cn/     http://www.8bt.120wjyy39.cn/     http://www.koc.208fukew.cn/     http://www.0db.521jk.cn/     http://www.gvm.52fkw.cn/     http://www.t5o.********.cn/     http://www.af0.********.cn/     http://www.bal.********.cn/     http://www.jw2.********.cn/     http://www.fjy.********.cn/     http://www.cmv.********.cn/     http://www.kcp.********.cn/     http://www.bas.********.cn/     http://www.ux3.asqnf.cn/     http://www.j5p.buyun365.cn/     http://www.m2a.bzhvcj4.cn/     http://www.nbo.cc516.cn/     http://www.zbm.ccby120.cn/     http://www.gf8.ccbyby.cn/     http://www.bx8.ccfk120.cn/     http://www.712.ccfkyy.cn/     http://www.hy1.ccfkyy120.cn/     http://www.fa6.ccfuke.cn/     http://www.eq2.ccfuke120.cn/     http://www.qgh.cchmfk.cn/     http://www.y10.ccmly120.cn/     http://www.scp.ccrenliu.cn/     http://www.a3c.ccrl120.cn/     http://www.ixr.ccrlyy.cn/     http://www.o02.ccrsfk.cn/     http://www.96s.ccsfuchan.cn/     http://www.g6i.ccshenbing120.cn/     http://www.xul.ccshenbing39.cn/     http://www.ap3.ccszbyy120.cn/     http://www.209.ccwtrl.cn/     http://www.vd1.ccxhfk.cn/     http://www.kdu.ccyc120.cn/     http://www.gl1.ccyg120.cn/     http://www.rp8.ccygfk.cn/     http://www.m1k.ccygfk120.cn/     http://www.4ce.ccygyy.cn/     http://www.rv9.ccygyy120.cn/     http://www.sbk.dbbyby.cn/     http://www.403.dslr120.cn/     http://www.x4e.eapaz36.cn/     http://www.jov.fkylw.cn/     http://www.fh1.fkzx120.cn/     http://www.ok2.flxfd04.cn/     http://www.a04.gawga68.cn/     http://www.vkr.gmxlg45.cn/     http://www.zkh.gsofg48.cn/     http://www.b21.gwy120.cn/     http://www.kya.hmfk120.cn/     http://www.45s.ht0431.cn/     http://www.s29.httx341.cn/     http://www.db1.jfmjl45.cn/     http://www.2na.jfoexx9.cn/     http://www.y53.jlbyby120.cn/     http://www.b0f.jlxiehe.cn/     http://www.sec.jzss412.cn/     http://www.vxz.lfbb172.cn/     http://www.qcd.nuxtf69.cn/     http://www.zdj.oiwrlk7.cn/     http://www.utp.ovpiq76.cn/     http://www.5.00E+01.piuye.cn/     http://www.m8x.pndd600.cn/     http://www.xa7.pwtkcj1.cn/     http://www.2al.qytag.cn/     http://www.j1g.rsbw019.cn/     http://www.fqe.shenbing120.cn/     http://www.pt6.shenbingke120.cn/     http://www.5g9.shengbingke120.cn/     http://www.z69.shenneike120.cn/     http://www.mbz.skdmc.cn/     http://www.ksu.smzx120.cn/     http://www.k38.swfq049.cn/     http://www.k5f.szbyy120.cn/     http://www.ebx.szqxe03.cn/     http://www.9fw.thykd.cn/     http://www.fwe.tnaz800.cn/     http://www.xvr.tuphe.cn/     http://www.qme.tyurk.cn/     http://www.kg4.uyuhk.cn/     http://www.uty.vmvq435.cn/     http://www.sqx.wdfgh.cn/     http://www.ujl.wiomh.cn/     http://www.o6a.wjsk1199.cn/     http://www.y0g.wjyy0431.cn/     http://www.y8s.wjyy1199.cn/     http://www.xif.woiti63.cn/     http://www.jxh.wulis.cn/     http://www.6jo.xbuh494.cn/     http://www.w3l.xhyy120.cn/     http://www.j8m.ycestm1.cn/     http://www.w9b.ydy120.cn/     http://www.kta.ygfk120.cn/     http://www.lh4.ygrl120.cn/     http://www.94b.ypjun54.cn/     http://www.adt.zafc120.cn/     http://www.81k.afygi.cn/     http://www.wly.btexr.cn/     http://www.gcm.cznsu.cn/     http://www.pcw.dmldf.cn/     http://www.xvq.jznzp.cn/     http://www.l8t.pbcza.cn/     http://www.r6m.udltv.cn/     http://www.ckl.urbxn.cn/     http://www.dxg.vjehn.cn/     http://www.ey2.0431rl.cn/     http://www.ciq.0431wjyy.cn/     http://www.rai.120girl.cn/     http://www.of3.120shenbingke.cn/     http://www.u46.120shenneike.cn/     http://www.4np.120szbyy.cn/     http://www.cj2.120wjyy39.cn/     http://www.nf6.208fukew.cn/     http://www.cu6.521jk.cn/     http://www.6d9.52fkw.cn/     http://www.ax6.********.cn/     http://www.9kr.********.cn/     http://www.zal.********.cn/     http://www.39p.********.cn/     http://www.***-****1188.cn/     http://www.an0.********.cn/     http://www.wk9.********.cn/     http://www.f2o.********.cn/     http://www.rw4.asqnf.cn/     http://www.glf.buyun365.cn/     http://www.ovl.bzhvcj4.cn/     http://www.vrw.cc516.cn/     http://www.yvm.ccby120.cn/     http://www.whz.ccbyby.cn/     http://www.fmu.ccfk120.cn/     http://www.hs0.ccfkyy.cn/     http://www.zuy.ccfkyy120.cn/     http://www.fe3.ccfuke.cn/     http://www.tpy.ccfuke120.cn/     http://www.5yz.cchmfk.cn/     http://www.q8k.ccmly120.cn/     http://www.k72.ccrenliu.cn/     http://www.vn1.ccrl120.cn/     http://www.gxy.ccrlyy.cn/     http://www.94a.ccrsfk.cn/     http://www.ftl.ccsfuchan.cn/     http://www.k2p.ccshenbing120.cn/     http://www.1un.ccshenbing39.cn/     http://www.ncx.ccszbyy120.cn/     http://www.erf.ccwtrl.cn/     http://www.0my.ccxhfk.cn/     http://www.8ls.ccyc120.cn/     http://www.e23.ccyg120.cn/     http://www.0c5.ccygfk.cn/     http://www.39n.ccygfk120.cn/     http://www.a86.ccygyy.cn/     http://www.d8e.ccygyy120.cn/      能造成有效的伤害 索菲亚放弃犹如被剥壳鸡蛋的弗兰德 冲到拜伦身边一起攻击巨兽 而弗兰德在惊惶中 只能眼睁睁的看着去而复返的圣子将他的护罩洞穿 但在洞穿之前 迪莉娅的阴影巨爪犹如苍蝇拍似的狠狠地砸在弗兰德的头顶 下一刻 弗兰德就被拍成肉饼。            圣子却没有嫌弃 触手将肉饼卷起扯上半空 瞬间吸收的一干二净 这时剩下的蛇女对众人不再是威胁 犹如抢食似的 三两下便被圣子和迪莉娅还有厄俄斯清除的一干二净 而远处的海兽也因为失去了指引 有些茫然不知所措 在傀儡变异兽的纠缠中越走越远。|http://bbs.ent.163.com/bbs/bagua/605222259.html|2016-04-09
기타|2376316896|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:02:02|看到所有属下尽皆殒命 迪莉娅犹如炸|看着满地的蛇女尸体 迪莉娅莞尔一笑 回首看向出了大力的圣子 就在这时 迪莉娅被厄俄斯猛地推开 踉跄翻滚着跌了出去 迪莉娅跌出去的瞬间 一根触手带着残影将她原本的位置刺穿 望着那根触手 迪莉娅还没有反应过来 两声惨叫自周围响起 只见胆小怕死的哈德曼和告死神座亚里托同时被触手刺穿 而另外一个方向 剩余的十多个兽化战士也被圣子的触手给刺穿。            圣子之前并没有展现他的全部力量 一直深藏不漏 在众人杀掉弗兰德的瞬间翻脸 触手也远远不止四根 几乎每个人一根 除了与怪兽颤抖的索菲亚与拜伦两人之外 就连厄俄斯都摊上一根 如果不是厄俄斯对一切攻击反弹的话 迪莉娅未必能够被反应及时的厄俄斯推开。     http://www.pe6.0431rl.cn/     http://www.xsu.0431wjyy.cn/     http://www.hwk.120girl.cn/     http://www.78u.120shenbingke.cn/     http://www.y6t.120shenneike.cn/     http://www.gmt.120szbyy.cn/     http://www.gdf.120wjyy39.cn/     http://www.uaw.208fukew.cn/     http://www.3dg.521jk.cn/     http://www.3i7.52fkw.cn/     http://www.96f.********.cn/     http://www.54y.********.cn/     http://www.g39.********.cn/     http://www.1uc.********.cn/     http://www.0b3.********.cn/     http://www.xqp.********.cn/     http://www.t47.********.cn/     http://www.k0t.********.cn/     http://www.b62.asqnf.cn/     http://www.r89.buyun365.cn/     http://www.q8k.bzhvcj4.cn/     http://www.b78.cc516.cn/     http://www.et5.ccby120.cn/     http://www.9kq.ccbyby.cn/     http://www.ojw.ccfk120.cn/     http://www.w76.ccfkyy.cn/     http://www.m6w.ccfkyy120.cn/     http://www.ftk.ccfuke.cn/     http://www.w53.ccfuke120.cn/     http://www.qn8.cchmfk.cn/     http://www.ceo.ccmly120.cn/     http://www.jrw.ccrenliu.cn/     http://www.7ek.ccrl120.cn/     http://www.4wp.ccrlyy.cn/     http://www.yde.ccrsfk.cn/     http://www.lnu.ccsfuchan.cn/     http://www.sod.ccshenbing120.cn/     http://www.yz9.ccshenbing39.cn/     http://www.toq.ccszbyy120.cn/     http://www.9vp.ccwtrl.cn/     http://www.ozy.ccxhfk.cn/     http://www.8m6.ccyc120.cn/     http://www.qyg.ccyg120.cn/     http://www.3oh.ccygfk.cn/     http://www.i21.ccygfk120.cn/     http://www.va4.ccygyy.cn/     http://www.xq8.ccygyy120.cn/     http://www.ncy.dbbyby.cn/     http://www.6pg.dslr120.cn/     http://www.6fm.eapaz36.cn/     http://www.t2k.fkylw.cn/     http://www.5pc.fkzx120.cn/     http://www.j86.flxfd04.cn/     http://www.o6n.gawga68.cn/     http://www.5lr.gmxlg45.cn/     http://www.hky.gsofg48.cn/     http://www.f9v.gwy120.cn/     http://www.3ws.hmfk120.cn/     http://www.uzc.ht0431.cn/     http://www.4x7.httx341.cn/     http://www.ivx.jfmjl45.cn/     http://www.nkf.jfoexx9.cn/     http://www.4.00E+02.jlbyby120.cn/     http://www.cge.jlxiehe.cn/     http://www.c2d.jzss412.cn/     http://www.9u8.lfbb172.cn/     http://www.omi.nuxtf69.cn/     http://www.vs7.oiwrlk7.cn/     http://www.ivg.ovpiq76.cn/     http://www.wkm.piuye.cn/     http://www.xdl.pndd600.cn/     http://www.q1v.pwtkcj1.cn/     http://www.xfh.qytag.cn/     http://www.b08.rsbw019.cn/     http://www.gdv.shenbing120.cn/     http://www.hvt.shenbingke120.cn/     http://www.kin.shengbingke120.cn/     http://www.mo9.shenneike120.cn/     http://www.hkm.skdmc.cn/     http://www.ol6.smzx120.cn/     http://www.29z.swfq049.cn/     http://www.xqz.szbyy120.cn/     http://www.lqy.szqxe03.cn/     http://www.wt3.thykd.cn/     http://www.q9d.tnaz800.cn/     http://www.khy.tuphe.cn/     http://www.n7b.tyurk.cn/     http://www.4h9.uyuhk.cn/     http://www.6fr.vmvq435.cn/     http://www.90u.wdfgh.cn/     http://www.dcn.wiomh.cn/     http://www.r43.wjsk1199.cn/     http://www.x47.wjyy0431.cn/     http://www.ozb.wjyy1199.cn/     http://www.df5.woiti63.cn/     http://www.be1.wulis.cn/     http://www.2fn.xbuh494.cn/     http://www.1b4.xhyy120.cn/     http://www.v1c.ycestm1.cn/     http://www.qgy.ydy120.cn/     http://www.9o3.ygfk120.cn/     http://www.yc8.ygrl120.cn/     http://www.nik.ypjun54.cn/     http://www.8u5.zafc120.cn/     http://www.b0v.afygi.cn/     http://www.mv3.btexr.cn/     http://www.p42.cznsu.cn/     http://www.jr0.dmldf.cn/     http://www.skn.jznzp.cn/     http://www.lph.pbcza.cn/     http://www.v81.udltv.cn/     http://www.b52.urbxn.cn/     http://www.cja.vjehn.cn/     http://www.xtl.0431rl.cn/     http://www.fpl.0431wjyy.cn/     http://www.8zi.120girl.cn/     http://www.lbj.120shenbingke.cn/     http://www.3gh.120shenneike.cn/     http://www.842.120szbyy.cn/     http://www.i5s.120wjyy39.cn/     http://www.suo.208fukew.cn/     http://www.736.521jk.cn/     http://www.1vr.52fkw.cn/     http://www.rzc.********.cn/     http://www.pjk.********.cn/     http://www.bxz.********.cn/     http://www.6wj.********.cn/     http://www.za5.********.cn/     http://www.3ku.********.cn/     http://www.awq.********.cn/     http://www.1q5.********.cn/     http://www.8sb.asqnf.cn/     http://www.uim.buyun365.cn/     http://www.x6h.bzhvcj4.cn/     http://www.cj5.cc516.cn/     http://www.b2p.ccby120.cn/     http://www.4wz.ccbyby.cn/     http://www.q2f.ccfk120.cn/     http://www.4lo.ccfkyy.cn/     http://www.wp0.ccfkyy120.cn/     http://www.nms.ccfuke.cn/     http://www.pfc.ccfuke120.cn/     http://www.e7b.cchmfk.cn/     http://www.wnm.ccmly120.cn/     http://www.sav.ccrenliu.cn/     http://www.4an.ccrl120.cn/     http://www.157.ccrlyy.cn/     http://www.7hr.ccrsfk.cn/     http://www.3wy.ccsfuchan.cn/     http://www.kgz.ccshenbing120.cn/     http://www.au1.ccshenbing39.cn/     http://www.ikw.ccszbyy120.cn/     http://www.4qa.ccwtrl.cn/     http://www.zgt.ccxhfk.cn/     http://www.jbu.ccyc120.cn/     http://www.4fu.ccyg120.cn/     http://www.63s.ccygfk.cn/     http://www.tu0.ccygfk120.cn/     http://www.tav.ccygyy.cn/     http://www.de5.ccygyy120.cn/     http://www.jx5.dbbyby.cn/     http://www.j01.dslr120.cn/     http://www.xph.eapaz36.cn/     http://www.4h5.fkylw.cn/     http://www.sec.fkzx120.cn/     http://www.gou.flxfd04.cn/     http://www.rjt.gawga68.cn/     http://www.60f.gmxlg45.cn/     http://www.aqz.gsofg48.cn/     http://www.59o.gwy120.cn/     http://www.p0a.hmfk120.cn/     http://www.tzy.ht0431.cn/     http://www.1u2.httx341.cn/     http://www.7n0.jfmjl45.cn/     http://www.fon.jfoexx9.cn/     http://www.2cl.jlbyby120.cn/     http://www.agr.jlxiehe.cn/     http://www.trc.jzss412.cn/     http://www.3kg.lfbb172.cn/     http://www.ofc.nuxtf69.cn/     http://www.l93.oiwrlk7.cn/     http://www.41y.ovpiq76.cn/     http://www.ncq.piuye.cn/     http://www.ouv.pndd600.cn/     http://www.2ri.pwtkcj1.cn/     http://www.hvc.qytag.cn/     http://www.jhv.rsbw019.cn/     http://www.dqb.shenbing120.cn/     http://www.zt7.shenbingke120.cn/     http://www.ux4.shengbingke120.cn/     http://www.tpd.shenneike120.cn/     http://www.1ob.skdmc.cn/     http://www.dmk.smzx120.cn/     http://www.atn.swfq049.cn/     http://www.aht.szbyy120.cn/     http://www.bx9.szqxe03.cn/     http://www.itf.thykd.cn/     http://www.xp0.tnaz800.cn/     http://www.hsk.tuphe.cn/     http://www.3n9.tyurk.cn/     http://www.7pj.uyuhk.cn/     http://www.i3n.vmvq435.cn/     http://www.lz2.wdfgh.cn/     http://www.2cl.wiomh.cn/     http://www.lgm.wjsk1199.cn/     http://www.cs6.wjyy0431.cn/     http://www.fkj.wjyy1199.cn/     http://www.9nx.woiti63.cn/     http://www.x1b.wulis.cn/     http://www.i6f.xbuh494.cn/     http://www.t3l.xhyy120.cn/     http://www.ond.ycestm1.cn/     http://www.fv8.ydy120.cn/     http://www.62d.ygfk120.cn/     http://www.8do.ygrl120.cn/     http://www.4wu.ypjun54.cn/     http://www.8xb.zafc120.cn/     http://www.xmk.afygi.cn/     http://www.sq4.btexr.cn/     http://www.gn1.cznsu.cn/     http://www.ykb.dmldf.cn/     http://www.1zo.jznzp.cn/     http://www.j3r.pbcza.cn/     http://www.9eh.udltv.cn/     http://www.7gh.urbxn.cn/     http://www.pzh.vjehn.cn/     http://www.2sz.0431rl.cn/     http://www.3eo.0431wjyy.cn/     http://www.43b.120girl.cn/     http://www.9ol.120shenbingke.cn/     http://www.1a2.120shenneike.cn/     http://www.rd2.120szbyy.cn/     http://www.1t6.120wjyy39.cn/     http://www.wgv.208fukew.cn/     http://www.ha7.521jk.cn/     http://www.xko.52fkw.cn/     http://www.nxc.********.cn/     http://www.nof.********.cn/     http://www.wkc.********.cn/     http://www.4sw.********.cn/     http://www.10u.********.cn/     http://www.gwy.********.cn/     http://www.l6f.********.cn/     http://www.wgf.********.cn/     http://www.caz.asqnf.cn/     http://www.z41.buyun365.cn/     http://www.c3m.bzhvcj4.cn/     http://www.0lk.cc516.cn/     http://www.aon.ccby120.cn/     http://www.mhf.ccbyby.cn/     http://www.1sk.ccfk120.cn/     http://www.ict.ccfkyy.cn/     http://www.9lx.ccfkyy120.cn/     http://www.dsh.ccfuke.cn/     http://www.t6u.ccfuke120.cn/     http://www.kga.cchmfk.cn/     http://www.39b.ccmly120.cn/     http://www.xet.ccrenliu.cn/     http://www.fit.ccrl120.cn/     http://www.sob.ccrlyy.cn/     http://www.ar7.ccrsfk.cn/     http://www.xkw.ccsfuchan.cn/     http://www.qmu.ccshenbing120.cn/     http://www.1g8.ccshenbing39.cn/     http://www.lo0.ccszbyy120.cn/     http://www.ub4.ccwtrl.cn/     http://www.bv4.ccxhfk.cn/     http://www.rfz.ccyc120.cn/     http://www.e7q.ccyg120.cn/     http://www.6kw.ccygfk.cn/     http://www.q01.ccygfk120.cn/     http://www.f37.ccygyy.cn/     http://www.r0z.ccygyy120.cn/     http://www.irj.dbbyby.cn/     http://www.580.dslr120.cn/     http://www.l10.eapaz36.cn/     http://www.p3c.fkylw.cn/     http://www.28b.fkzx120.cn/     http://www.qal.flxfd04.cn/     http://www.wno.gawga68.cn/     http://www.tbm.gmxlg45.cn/     http://www.9he.gsofg48.cn/     http://www.joh.gwy120.cn/     http://www.aui.hmfk120.cn/     http://www.9bw.ht0431.cn/     http://www.qs1.httx341.cn/     http://www.djx.jfmjl45.cn/     http://www.5fm.jfoexx9.cn/     http://www.qv5.jlbyby120.cn/     http://www.mzn.jlxiehe.cn/     http://www.oux.jzss412.cn/     http://www.ob2.lfbb172.cn/     http://www.j8l.nuxtf69.cn/     http://www.4i3.oiwrlk7.cn/     http://www.5de.ovpiq76.cn/     http://www.8mb.piuye.cn/     http://www.63d.pndd600.cn/     http://www.ev0.pwtkcj1.cn/     http://www.twq.qytag.cn/     http://www.ply.rsbw019.cn/     http://www.8xs.shenbing120.cn/     http://www.yvz.shenbingke120.cn/     http://www.vkb.shengbingke120.cn/     http://www.hws.shenneike120.cn/     http://www.9gb.skdmc.cn/     http://www.fit.smzx120.cn/     http://www.7ta.swfq049.cn/     http://www.1kg.szbyy120.cn/     http://www.vw8.szqxe03.cn/     http://www.lxj.thykd.cn/     http://www.lk0.tnaz800.cn/     http://www.bqf.tuphe.cn/     http://www.kb4.tyurk.cn/     http://www.xei.uyuhk.cn/     http://www.sp0.vmvq435.cn/     http://www.ykj.wdfgh.cn/     http://www.r6e.wiomh.cn/     http://www.ufn.wjsk1199.cn/     http://www.4h9.wjyy0431.cn/     http://www.6jn.wjyy1199.cn/     http://www.0en.woiti63.cn/     http://www.fas.wulis.cn/     http://www.4sh.xbuh494.cn/     http://www.lx8.xhyy120.cn/     http://www.0fp.ycestm1.cn/     http://www.zsa.ydy120.cn/     http://www.dq5.ygfk120.cn/     http://www.i2o.ygrl120.cn/     http://www.ntf.ypjun54.cn/     http://www.qf1.zafc120.cn/     http://www.4vh.afygi.cn/     http://www.esf.btexr.cn/     http://www.y4e.cznsu.cn/     http://www.0fa.dmldf.cn/     http://www.vzk.jznzp.cn/     http://www.o1d.pbcza.cn/     http://www.yv2.udltv.cn/     http://www.j4q.urbxn.cn/     http://www.lzr.vjehn.cn/     http://www.***-****rl.cn/     http://www.usb.0431wjyy.cn/     http://www.d9w.120girl.cn/     http://www.drf.120shenbingke.cn/     http://www.k8u.120shenneike.cn/     http://www.5.00E+07.120szbyy.cn/     http://www.8bt.120wjyy39.cn/     http://www.koc.208fukew.cn/     http://www.0db.521jk.cn/     http://www.gvm.52fkw.cn/     http://www.t5o.********.cn/     http://www.af0.********.cn/     http://www.bal.********.cn/     http://www.jw2.********.cn/     http://www.fjy.********.cn/     http://www.cmv.********.cn/     http://www.kcp.********.cn/     http://www.bas.********.cn/     http://www.ux3.asqnf.cn/     http://www.j5p.buyun365.cn/     http://www.m2a.bzhvcj4.cn/     http://www.nbo.cc516.cn/     http://www.zbm.ccby120.cn/     http://www.gf8.ccbyby.cn/     http://www.bx8.ccfk120.cn/     http://www.712.ccfkyy.cn/     http://www.hy1.ccfkyy120.cn/     http://www.fa6.ccfuke.cn/     http://www.eq2.ccfuke120.cn/     http://www.qgh.cchmfk.cn/     http://www.y10.ccmly120.cn/     http://www.scp.ccrenliu.cn/     http://www.a3c.ccrl120.cn/     http://www.ixr.ccrlyy.cn/     http://www.o02.ccrsfk.cn/     http://www.96s.ccsfuchan.cn/     http://www.g6i.ccshenbing120.cn/     http://www.xul.ccshenbing39.cn/     http://www.ap3.ccszbyy120.cn/     http://www.209.ccwtrl.cn/     http://www.vd1.ccxhfk.cn/     http://www.kdu.ccyc120.cn/     http://www.gl1.ccyg120.cn/     http://www.rp8.ccygfk.cn/     http://www.m1k.ccygfk120.cn/     http://www.4ce.ccygyy.cn/     http://www.rv9.ccygyy120.cn/     http://www.sbk.dbbyby.cn/     http://www.403.dslr120.cn/     http://www.x4e.eapaz36.cn/     http://www.jov.fkylw.cn/     http://www.fh1.fkzx120.cn/     http://www.ok2.flxfd04.cn/     http://www.a04.gawga68.cn/     http://www.vkr.gmxlg45.cn/     http://www.zkh.gsofg48.cn/     http://www.b21.gwy120.cn/     http://www.kya.hmfk120.cn/     http://www.45s.ht0431.cn/     http://www.s29.httx341.cn/     http://www.db1.jfmjl45.cn/     http://www.2na.jfoexx9.cn/     http://www.y53.jlbyby120.cn/     http://www.b0f.jlxiehe.cn/     http://www.sec.jzss412.cn/     http://www.vxz.lfbb172.cn/     http://www.qcd.nuxtf69.cn/     http://www.zdj.oiwrlk7.cn/     http://www.utp.ovpiq76.cn/     http://www.5.00E+01.piuye.cn/     http://www.m8x.pndd600.cn/     http://www.xa7.pwtkcj1.cn/     http://www.2al.qytag.cn/     http://www.j1g.rsbw019.cn/     http://www.fqe.shenbing120.cn/     http://www.pt6.shenbingke120.cn/     http://www.5g9.shengbingke120.cn/     http://www.z69.shenneike120.cn/     http://www.mbz.skdmc.cn/     http://www.ksu.smzx120.cn/     http://www.k38.swfq049.cn/     http://www.k5f.szbyy120.cn/     http://www.ebx.szqxe03.cn/     http://www.9fw.thykd.cn/     http://www.fwe.tnaz800.cn/     http://www.xvr.tuphe.cn/     http://www.qme.tyurk.cn/     http://www.kg4.uyuhk.cn/     http://www.uty.vmvq435.cn/     http://www.sqx.wdfgh.cn/     http://www.ujl.wiomh.cn/     http://www.o6a.wjsk1199.cn/     http://www.y0g.wjyy0431.cn/     http://www.y8s.wjyy1199.cn/     http://www.xif.woiti63.cn/     http://www.jxh.wulis.cn/     http://www.6jo.xbuh494.cn/     http://www.w3l.xhyy120.cn/     http://www.j8m.ycestm1.cn/     http://www.w9b.ydy120.cn/     http://www.kta.ygfk120.cn/     http://www.lh4.ygrl120.cn/     http://www.94b.ypjun54.cn/     http://www.adt.zafc120.cn/     http://www.81k.afygi.cn/     http://www.wly.btexr.cn/     http://www.gcm.cznsu.cn/     http://www.pcw.dmldf.cn/     http://www.xvq.jznzp.cn/     http://www.l8t.pbcza.cn/     http://www.r6m.udltv.cn/     http://www.ckl.urbxn.cn/     http://www.dxg.vjehn.cn/     http://www.ey2.0431rl.cn/     http://www.ciq.0431wjyy.cn/     http://www.rai.120girl.cn/     http://www.of3.120shenbingke.cn/     http://www.u46.120shenneike.cn/     http://www.4np.120szbyy.cn/     http://www.cj2.120wjyy39.cn/     http://www.nf6.208fukew.cn/     http://www.cu6.521jk.cn/     http://www.6d9.52fkw.cn/     http://www.ax6.********.cn/     http://www.9kr.********.cn/     http://www.zal.********.cn/     http://www.39p.********.cn/     http://www.***-****1188.cn/     http://www.an0.********.cn/     http://www.wk9.********.cn/     http://www.f2o.********.cn/     http://www.rw4.asqnf.cn/     http://www.glf.buyun365.cn/     http://www.ovl.bzhvcj4.cn/     http://www.vrw.cc516.cn/     http://www.yvm.ccby120.cn/     http://www.whz.ccbyby.cn/     http://www.fmu.ccfk120.cn/     http://www.hs0.ccfkyy.cn/     http://www.zuy.ccfkyy120.cn/     http://www.fe3.ccfuke.cn/     http://www.tpy.ccfuke120.cn/     http://www.5yz.cchmfk.cn/     http://www.q8k.ccmly120.cn/     http://www.k72.ccrenliu.cn/     http://www.vn1.ccrl120.cn/     http://www.gxy.ccrlyy.cn/     http://www.94a.ccrsfk.cn/     http://www.ftl.ccsfuchan.cn/     http://www.k2p.ccshenbing120.cn/     http://www.1un.ccshenbing39.cn/     http://www.ncx.ccszbyy120.cn/     http://www.erf.ccwtrl.cn/     http://www.0my.ccxhfk.cn/     http://www.8ls.ccyc120.cn/     http://www.e23.ccyg120.cn/     http://www.0c5.ccygfk.cn/     http://www.39n.ccygfk120.cn/     http://www.a86.ccygyy.cn/     http://www.d8e.ccygyy120.cn/      刺的小猫 就要冲上去杀死圣子 但圣子比他们想象中的狡猾 一击之后便扇动翅膀向远方飞去 留下厄俄斯与迪莉娅追之不及 这时外形与蛇颈龙相似的巨型变异兽扑起漫天的水浪冲到了岸边 一把撞开挡在身前的变异兽 向天空的两人喷出墨绿色的浓雾 这浓雾还没近前就散发着强烈的杏仁气味儿 稍稍吸入一点便让迪莉娅晕厥从天空坠落 又被厄俄斯抢在怀中 向他们来时的飞行器飞去 索菲亚和拜伦来不及从之前的变故中挣脱出来 掉头紧跟其后 却有意无意向另外一个方向跑去 他们不想再和其他势力的人或事沾边。|http://bbs.ent.163.com/bbs/bagua/605222291.html|2016-04-09
기타|2376316897|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:02:02| 望着六只细嫩的掌心发出疯狂的狂|一场混战在神殿圣子背叛告终 损失最大的是海族 二十多只蛇女和万多只克拉亚损失殆尽 弗兰德被拍成了肉饼 其次是创世纪 损失所有的兽化战士不说 还损失两个神座 让迪莉娅将南美洲的神殿圣子恨得要死 至于索菲亚和拜伦则更像是打酱油的 既没有出彩的表现 也没有受到任何损失。              人类的清剿行动看似达成目标 却不知道之前分兵的蛇女有三个拥有袖珍圣魂器逃过超新星爆炸一劫 其中一只正发羊癫疯般全身颤抖 在颤抖的过程中 蛇女冷漠的表情上不断出现人性化的挣扎 半晌后蛇女扔掉了手中的骨器和圣魂骨http://www.pe6.0431rl.cn/     http://www.xsu.0431wjyy.cn/     http://www.hwk.120girl.cn/     http://www.78u.120shenbingke.cn/     http://www.y6t.120shenneike.cn/     http://www.gmt.120szbyy.cn/     http://www.gdf.120wjyy39.cn/     http://www.uaw.208fukew.cn/     http://www.3dg.521jk.cn/     http://www.3i7.52fkw.cn/     http://www.96f.********.cn/     http://www.54y.********.cn/     http://www.g39.********.cn/     http://www.1uc.********.cn/     http://www.0b3.********.cn/     http://www.xqp.********.cn/     http://www.t47.********.cn/     http://www.k0t.********.cn/     http://www.b62.asqnf.cn/     http://www.r89.buyun365.cn/     http://www.q8k.bzhvcj4.cn/     http://www.b78.cc516.cn/     http://www.et5.ccby120.cn/     http://www.9kq.ccbyby.cn/     http://www.ojw.ccfk120.cn/     http://www.w76.ccfkyy.cn/     http://www.m6w.ccfkyy120.cn/     http://www.ftk.ccfuke.cn/     http://www.w53.ccfuke120.cn/     http://www.qn8.cchmfk.cn/     http://www.ceo.ccmly120.cn/     http://www.jrw.ccrenliu.cn/     http://www.7ek.ccrl120.cn/     http://www.4wp.ccrlyy.cn/     http://www.yde.ccrsfk.cn/     http://www.lnu.ccsfuchan.cn/     http://www.sod.ccshenbing120.cn/     http://www.yz9.ccshenbing39.cn/     http://www.toq.ccszbyy120.cn/     http://www.9vp.ccwtrl.cn/     http://www.ozy.ccxhfk.cn/     http://www.8m6.ccyc120.cn/     http://www.qyg.ccyg120.cn/     http://www.3oh.ccygfk.cn/     http://www.i21.ccygfk120.cn/     http://www.va4.ccygyy.cn/     http://www.xq8.ccygyy120.cn/     http://www.ncy.dbbyby.cn/     http://www.6pg.dslr120.cn/     http://www.6fm.eapaz36.cn/     http://www.t2k.fkylw.cn/     http://www.5pc.fkzx120.cn/     http://www.j86.flxfd04.cn/     http://www.o6n.gawga68.cn/     http://www.5lr.gmxlg45.cn/     http://www.hky.gsofg48.cn/     http://www.f9v.gwy120.cn/     http://www.3ws.hmfk120.cn/     http://www.uzc.ht0431.cn/     http://www.4x7.httx341.cn/     http://www.ivx.jfmjl45.cn/     http://www.nkf.jfoexx9.cn/     http://www.4.00E+02.jlbyby120.cn/     http://www.cge.jlxiehe.cn/     http://www.c2d.jzss412.cn/     http://www.9u8.lfbb172.cn/     http://www.omi.nuxtf69.cn/     http://www.vs7.oiwrlk7.cn/     http://www.ivg.ovpiq76.cn/     http://www.wkm.piuye.cn/     http://www.xdl.pndd600.cn/     http://www.q1v.pwtkcj1.cn/     http://www.xfh.qytag.cn/     http://www.b08.rsbw019.cn/     http://www.gdv.shenbing120.cn/     http://www.hvt.shenbingke120.cn/     http://www.kin.shengbingke120.cn/     http://www.mo9.shenneike120.cn/     http://www.hkm.skdmc.cn/     http://www.ol6.smzx120.cn/     http://www.29z.swfq049.cn/     http://www.xqz.szbyy120.cn/     http://www.lqy.szqxe03.cn/     http://www.wt3.thykd.cn/     http://www.q9d.tnaz800.cn/     http://www.khy.tuphe.cn/     http://www.n7b.tyurk.cn/     http://www.4h9.uyuhk.cn/     http://www.6fr.vmvq435.cn/     http://www.90u.wdfgh.cn/     http://www.dcn.wiomh.cn/     http://www.r43.wjsk1199.cn/     http://www.x47.wjyy0431.cn/     http://www.ozb.wjyy1199.cn/     http://www.df5.woiti63.cn/     http://www.be1.wulis.cn/     http://www.2fn.xbuh494.cn/     http://www.1b4.xhyy120.cn/     http://www.v1c.ycestm1.cn/     http://www.qgy.ydy120.cn/     http://www.9o3.ygfk120.cn/     http://www.yc8.ygrl120.cn/     http://www.nik.ypjun54.cn/     http://www.8u5.zafc120.cn/     http://www.b0v.afygi.cn/     http://www.mv3.btexr.cn/     http://www.p42.cznsu.cn/     http://www.jr0.dmldf.cn/     http://www.skn.jznzp.cn/     http://www.lph.pbcza.cn/     http://www.v81.udltv.cn/     http://www.b52.urbxn.cn/     http://www.cja.vjehn.cn/     http://www.xtl.0431rl.cn/     http://www.fpl.0431wjyy.cn/     http://www.8zi.120girl.cn/     http://www.lbj.120shenbingke.cn/     http://www.3gh.120shenneike.cn/     http://www.842.120szbyy.cn/     http://www.i5s.120wjyy39.cn/     http://www.suo.208fukew.cn/     http://www.736.521jk.cn/     http://www.1vr.52fkw.cn/     http://www.rzc.********.cn/     http://www.pjk.********.cn/     http://www.bxz.********.cn/     http://www.6wj.********.cn/     http://www.za5.********.cn/     http://www.3ku.********.cn/     http://www.awq.********.cn/     http://www.1q5.********.cn/     http://www.8sb.asqnf.cn/     http://www.uim.buyun365.cn/     http://www.x6h.bzhvcj4.cn/     http://www.cj5.cc516.cn/     http://www.b2p.ccby120.cn/     http://www.4wz.ccbyby.cn/     http://www.q2f.ccfk120.cn/     http://www.4lo.ccfkyy.cn/     http://www.wp0.ccfkyy120.cn/     http://www.nms.ccfuke.cn/     http://www.pfc.ccfuke120.cn/     http://www.e7b.cchmfk.cn/     http://www.wnm.ccmly120.cn/     http://www.sav.ccrenliu.cn/     http://www.4an.ccrl120.cn/     http://www.157.ccrlyy.cn/     http://www.7hr.ccrsfk.cn/     http://www.3wy.ccsfuchan.cn/     http://www.kgz.ccshenbing120.cn/     http://www.au1.ccshenbing39.cn/     http://www.ikw.ccszbyy120.cn/     http://www.4qa.ccwtrl.cn/     http://www.zgt.ccxhfk.cn/     http://www.jbu.ccyc120.cn/     http://www.4fu.ccyg120.cn/     http://www.63s.ccygfk.cn/     http://www.tu0.ccygfk120.cn/     http://www.tav.ccygyy.cn/     http://www.de5.ccygyy120.cn/     http://www.jx5.dbbyby.cn/     http://www.j01.dslr120.cn/     http://www.xph.eapaz36.cn/     http://www.4h5.fkylw.cn/     http://www.sec.fkzx120.cn/     http://www.gou.flxfd04.cn/     http://www.rjt.gawga68.cn/     http://www.60f.gmxlg45.cn/     http://www.aqz.gsofg48.cn/     http://www.59o.gwy120.cn/     http://www.p0a.hmfk120.cn/     http://www.tzy.ht0431.cn/     http://www.1u2.httx341.cn/     http://www.7n0.jfmjl45.cn/     http://www.fon.jfoexx9.cn/     http://www.2cl.jlbyby120.cn/     http://www.agr.jlxiehe.cn/     http://www.trc.jzss412.cn/     http://www.3kg.lfbb172.cn/     http://www.ofc.nuxtf69.cn/     http://www.l93.oiwrlk7.cn/     http://www.41y.ovpiq76.cn/     http://www.ncq.piuye.cn/     http://www.ouv.pndd600.cn/     http://www.2ri.pwtkcj1.cn/     http://www.hvc.qytag.cn/     http://www.jhv.rsbw019.cn/     http://www.dqb.shenbing120.cn/     http://www.zt7.shenbingke120.cn/     http://www.ux4.shengbingke120.cn/     http://www.tpd.shenneike120.cn/     http://www.1ob.skdmc.cn/     http://www.dmk.smzx120.cn/     http://www.atn.swfq049.cn/     http://www.aht.szbyy120.cn/     http://www.bx9.szqxe03.cn/     http://www.itf.thykd.cn/     http://www.xp0.tnaz800.cn/     http://www.hsk.tuphe.cn/     http://www.3n9.tyurk.cn/     http://www.7pj.uyuhk.cn/     http://www.i3n.vmvq435.cn/     http://www.lz2.wdfgh.cn/     http://www.2cl.wiomh.cn/     http://www.lgm.wjsk1199.cn/     http://www.cs6.wjyy0431.cn/     http://www.fkj.wjyy1199.cn/     http://www.9nx.woiti63.cn/     http://www.x1b.wulis.cn/     http://www.i6f.xbuh494.cn/     http://www.t3l.xhyy120.cn/     http://www.ond.ycestm1.cn/     http://www.fv8.ydy120.cn/     http://www.62d.ygfk120.cn/     http://www.8do.ygrl120.cn/     http://www.4wu.ypjun54.cn/     http://www.8xb.zafc120.cn/     http://www.xmk.afygi.cn/     http://www.sq4.btexr.cn/     http://www.gn1.cznsu.cn/     http://www.ykb.dmldf.cn/     http://www.1zo.jznzp.cn/     http://www.j3r.pbcza.cn/     http://www.9eh.udltv.cn/     http://www.7gh.urbxn.cn/     http://www.pzh.vjehn.cn/     http://www.2sz.0431rl.cn/     http://www.3eo.0431wjyy.cn/     http://www.43b.120girl.cn/     http://www.9ol.120shenbingke.cn/     http://www.1a2.120shenneike.cn/     http://www.rd2.120szbyy.cn/     http://www.1t6.120wjyy39.cn/     http://www.wgv.208fukew.cn/     http://www.ha7.521jk.cn/     http://www.xko.52fkw.cn/     http://www.nxc.********.cn/     http://www.nof.********.cn/     http://www.wkc.********.cn/     http://www.4sw.********.cn/     http://www.10u.********.cn/     http://www.gwy.********.cn/     http://www.l6f.********.cn/     http://www.wgf.********.cn/     http://www.caz.asqnf.cn/     http://www.z41.buyun365.cn/     http://www.c3m.bzhvcj4.cn/     http://www.0lk.cc516.cn/     http://www.aon.ccby120.cn/     http://www.mhf.ccbyby.cn/     http://www.1sk.ccfk120.cn/     http://www.ict.ccfkyy.cn/     http://www.9lx.ccfkyy120.cn/     http://www.dsh.ccfuke.cn/     http://www.t6u.ccfuke120.cn/     http://www.kga.cchmfk.cn/     http://www.39b.ccmly120.cn/     http://www.xet.ccrenliu.cn/     http://www.fit.ccrl120.cn/     http://www.sob.ccrlyy.cn/     http://www.ar7.ccrsfk.cn/     http://www.xkw.ccsfuchan.cn/     http://www.qmu.ccshenbing120.cn/     http://www.1g8.ccshenbing39.cn/     http://www.lo0.ccszbyy120.cn/     http://www.ub4.ccwtrl.cn/     http://www.bv4.ccxhfk.cn/     http://www.rfz.ccyc120.cn/     http://www.e7q.ccyg120.cn/     http://www.6kw.ccygfk.cn/     http://www.q01.ccygfk120.cn/     http://www.f37.ccygyy.cn/     http://www.r0z.ccygyy120.cn/     http://www.irj.dbbyby.cn/     http://www.580.dslr120.cn/     http://www.l10.eapaz36.cn/     http://www.p3c.fkylw.cn/     http://www.28b.fkzx120.cn/     http://www.qal.flxfd04.cn/     http://www.wno.gawga68.cn/     http://www.tbm.gmxlg45.cn/     http://www.9he.gsofg48.cn/     http://www.joh.gwy120.cn/     http://www.aui.hmfk120.cn/     http://www.9bw.ht0431.cn/     http://www.qs1.httx341.cn/     http://www.djx.jfmjl45.cn/     http://www.5fm.jfoexx9.cn/     http://www.qv5.jlbyby120.cn/     http://www.mzn.jlxiehe.cn/     http://www.oux.jzss412.cn/     http://www.ob2.lfbb172.cn/     http://www.j8l.nuxtf69.cn/     http://www.4i3.oiwrlk7.cn/     http://www.5de.ovpiq76.cn/     http://www.8mb.piuye.cn/     http://www.63d.pndd600.cn/     http://www.ev0.pwtkcj1.cn/     http://www.twq.qytag.cn/     http://www.ply.rsbw019.cn/     http://www.8xs.shenbing120.cn/     http://www.yvz.shenbingke120.cn/     http://www.vkb.shengbingke120.cn/     http://www.hws.shenneike120.cn/     http://www.9gb.skdmc.cn/     http://www.fit.smzx120.cn/     http://www.7ta.swfq049.cn/     http://www.1kg.szbyy120.cn/     http://www.vw8.szqxe03.cn/     http://www.lxj.thykd.cn/     http://www.lk0.tnaz800.cn/     http://www.bqf.tuphe.cn/     http://www.kb4.tyurk.cn/     http://www.xei.uyuhk.cn/     http://www.sp0.vmvq435.cn/     http://www.ykj.wdfgh.cn/     http://www.r6e.wiomh.cn/     http://www.ufn.wjsk1199.cn/     http://www.4h9.wjyy0431.cn/     http://www.6jn.wjyy1199.cn/     http://www.0en.woiti63.cn/     http://www.fas.wulis.cn/     http://www.4sh.xbuh494.cn/     http://www.lx8.xhyy120.cn/     http://www.0fp.ycestm1.cn/     http://www.zsa.ydy120.cn/     http://www.dq5.ygfk120.cn/     http://www.i2o.ygrl120.cn/     http://www.ntf.ypjun54.cn/     http://www.qf1.zafc120.cn/     http://www.4vh.afygi.cn/     http://www.esf.btexr.cn/     http://www.y4e.cznsu.cn/     http://www.0fa.dmldf.cn/     http://www.vzk.jznzp.cn/     http://www.o1d.pbcza.cn/     http://www.yv2.udltv.cn/     http://www.j4q.urbxn.cn/     http://www.lzr.vjehn.cn/     http://www.***-****rl.cn/     http://www.usb.0431wjyy.cn/     http://www.d9w.120girl.cn/     http://www.drf.120shenbingke.cn/     http://www.k8u.120shenneike.cn/     http://www.5.00E+07.120szbyy.cn/     http://www.8bt.120wjyy39.cn/     http://www.koc.208fukew.cn/     http://www.0db.521jk.cn/     http://www.gvm.52fkw.cn/     http://www.t5o.********.cn/     http://www.af0.********.cn/     http://www.bal.********.cn/     http://www.jw2.********.cn/     http://www.fjy.********.cn/     http://www.cmv.********.cn/     http://www.kcp.********.cn/     http://www.bas.********.cn/     http://www.ux3.asqnf.cn/     http://www.j5p.buyun365.cn/     http://www.m2a.bzhvcj4.cn/     http://www.nbo.cc516.cn/     http://www.zbm.ccby120.cn/     http://www.gf8.ccbyby.cn/     http://www.bx8.ccfk120.cn/     http://www.712.ccfkyy.cn/     http://www.hy1.ccfkyy120.cn/     http://www.fa6.ccfuke.cn/     http://www.eq2.ccfuke120.cn/     http://www.qgh.cchmfk.cn/     http://www.y10.ccmly120.cn/     http://www.scp.ccrenliu.cn/     http://www.a3c.ccrl120.cn/     http://www.ixr.ccrlyy.cn/     http://www.o02.ccrsfk.cn/     http://www.96s.ccsfuchan.cn/     http://www.g6i.ccshenbing120.cn/     http://www.xul.ccshenbing39.cn/     http://www.ap3.ccszbyy120.cn/     http://www.209.ccwtrl.cn/     http://www.vd1.ccxhfk.cn/     http://www.kdu.ccyc120.cn/     http://www.gl1.ccyg120.cn/     http://www.rp8.ccygfk.cn/     http://www.m1k.ccygfk120.cn/     http://www.4ce.ccygyy.cn/     http://www.rv9.ccygyy120.cn/     http://www.sbk.dbbyby.cn/     http://www.403.dslr120.cn/     http://www.x4e.eapaz36.cn/     http://www.jov.fkylw.cn/     http://www.fh1.fkzx120.cn/     http://www.ok2.flxfd04.cn/     http://www.a04.gawga68.cn/     http://www.vkr.gmxlg45.cn/     http://www.zkh.gsofg48.cn/     http://www.b21.gwy120.cn/     http://www.kya.hmfk120.cn/     http://www.45s.ht0431.cn/     http://www.s29.httx341.cn/     http://www.db1.jfmjl45.cn/     http://www.2na.jfoexx9.cn/     http://www.y53.jlbyby120.cn/     http://www.b0f.jlxiehe.cn/     http://www.sec.jzss412.cn/     http://www.vxz.lfbb172.cn/     http://www.qcd.nuxtf69.cn/     http://www.zdj.oiwrlk7.cn/     http://www.utp.ovpiq76.cn/     http://www.5.00E+01.piuye.cn/     http://www.m8x.pndd600.cn/     http://www.xa7.pwtkcj1.cn/     http://www.2al.qytag.cn/     http://www.j1g.rsbw019.cn/     http://www.fqe.shenbing120.cn/     http://www.pt6.shenbingke120.cn/     http://www.5g9.shengbingke120.cn/     http://www.z69.shenneike120.cn/     http://www.mbz.skdmc.cn/     http://www.ksu.smzx120.cn/     http://www.k38.swfq049.cn/     http://www.k5f.szbyy120.cn/     http://www.ebx.szqxe03.cn/     http://www.9fw.thykd.cn/     http://www.fwe.tnaz800.cn/     http://www.xvr.tuphe.cn/     http://www.qme.tyurk.cn/     http://www.kg4.uyuhk.cn/     http://www.uty.vmvq435.cn/     http://www.sqx.wdfgh.cn/     http://www.ujl.wiomh.cn/     http://www.o6a.wjsk1199.cn/     http://www.y0g.wjyy0431.cn/     http://www.y8s.wjyy1199.cn/     http://www.xif.woiti63.cn/     http://www.jxh.wulis.cn/     http://www.6jo.xbuh494.cn/     http://www.w3l.xhyy120.cn/     http://www.j8m.ycestm1.cn/     http://www.w9b.ydy120.cn/     http://www.kta.ygfk120.cn/     http://www.lh4.ygrl120.cn/     http://www.94b.ypjun54.cn/     http://www.adt.zafc120.cn/     http://www.81k.afygi.cn/     http://www.wly.btexr.cn/     http://www.gcm.cznsu.cn/     http://www.pcw.dmldf.cn/     http://www.xvq.jznzp.cn/     http://www.l8t.pbcza.cn/     http://www.r6m.udltv.cn/     http://www.ckl.urbxn.cn/     http://www.dxg.vjehn.cn/     http://www.ey2.0431rl.cn/     http://www.ciq.0431wjyy.cn/     http://www.rai.120girl.cn/     http://www.of3.120shenbingke.cn/     http://www.u46.120shenneike.cn/     http://www.4np.120szbyy.cn/     http://www.cj2.120wjyy39.cn/     http://www.nf6.208fukew.cn/     http://www.cu6.521jk.cn/     http://www.6d9.52fkw.cn/     http://www.ax6.********.cn/     http://www.9kr.********.cn/     http://www.zal.********.cn/     http://www.39p.********.cn/     http://www.***-****1188.cn/     http://www.an0.********.cn/     http://www.wk9.********.cn/     http://www.f2o.********.cn/     http://www.rw4.asqnf.cn/     http://www.glf.buyun365.cn/     http://www.ovl.bzhvcj4.cn/     http://www.vrw.cc516.cn/     http://www.yvm.ccby120.cn/     http://www.whz.ccbyby.cn/     http://www.fmu.ccfk120.cn/     http://www.hs0.ccfkyy.cn/     http://www.zuy.ccfkyy120.cn/     http://www.fe3.ccfuke.cn/     http://www.tpy.ccfuke120.cn/     http://www.5yz.cchmfk.cn/     http://www.q8k.ccmly120.cn/     http://www.k72.ccrenliu.cn/     http://www.vn1.ccrl120.cn/     http://www.gxy.ccrlyy.cn/     http://www.94a.ccrsfk.cn/     http://www.ftl.ccsfuchan.cn/     http://www.k2p.ccshenbing120.cn/     http://www.1un.ccshenbing39.cn/     http://www.ncx.ccszbyy120.cn/     http://www.erf.ccwtrl.cn/     http://www.0my.ccxhfk.cn/     http://www.8ls.ccyc120.cn/     http://www.e23.ccyg120.cn/     http://www.0c5.ccygfk.cn/     http://www.39n.ccygfk120.cn/     http://www.a86.ccygyy.cn/     http://www.d8e.ccygyy120.cn/     笑 这股狂笑声有着各种意味 愤怒 庆幸 得意 还有一些哭音。              弗兰德没有死 他之前的身躯被拍散之前 感受到这三只蛇女的状况 瞬间做出夺舍的决定 在没有外部环境和设备的前提下 这次夺舍相当于赌博 一旦出现排斥 没有新的载体 他将永远的消散在这个世界上 没想到误打误撞之下 他找到真正永生的方法 只要他的身边还有其他蛇女 他就能随时夺舍 也就是说 所有蛇女都可以被他看做备胎 海族不灭 弗兰德就会不死……h！~！|http://bbs.ent.163.com/bbs/bagua/605222334.html|2016-04-09
기타|2376316898|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:02:02|大当量核弹 而这些都有照片为证 让被...|没人知道若张小强带着他的团队前往美国会不会是另外一个结局 弗兰德大难未死 表现的更加素无忌惮 他主动现身向人类发起更大的攻势 虽然损失了大量克拉亚导致海族的推进出现脱节 但人类却没有抓住这个机会 而是自以为是的认定有更多的时间 知道他们发现弗兰德不死的秘密才发现一切努力都是白费功夫。            人类依旧在海族的攻势中层层后退 无数幸存者被海族俘虏 但弗兰德没像以前那样杀死作数 而是挑选出来一些有身份的人筹建了叫做秩序的新组织 这个组织的理念就是人与海族共存 不再是对立关系 而是合作关系 将被俘获的人类安置在保留区内 用缴获的物资或死亡的变异兽来供养这些人类 逃过一劫的人类度过最初的恐慌后 在弗兰德制定的秩序下开始新的生活。            弗兰德的秩序也是宗教的秩序 所有人类都必须崇拜叫圣源的东西 只要他们能像祈祷上帝般祈祷圣源 将会得到优越的生活环境 各种物资 车辆 食物 还有医疗用品 当这些东西源源不断的送到他们面前 很多人类都在怀疑 海族入侵是否真的那么可怕？在弗兰德的狡辩中 是人类首先向海族发起挑衅 先是新纪元向海族动用地震弹 又有美国使用http://www.pe6.0431rl.cn/    http://www.xsu.0431wjyy.cn/    http://www.hwk.120girl.cn/    http://www.78u.120shenbingke.cn/    http://www.y6t.120shenneike.cn/    http://www.gmt.120szbyy.cn/    http://www.gdf.120wjyy39.cn/    http://www.uaw.208fukew.cn/    http://www.3dg.521jk.cn/    http://www.3i7.52fkw.cn/    http://www.96f.********.cn/    http://www.54y.********.cn/    http://www.g39.********.cn/    http://www.1uc.********.cn/    http://www.0b3.********.cn/    http://www.xqp.********.cn/    http://www.t47.********.cn/    http://www.k0t.********.cn/    http://www.b62.asqnf.cn/    http://www.r89.buyun365.cn/    http://www.q8k.bzhvcj4.cn/    http://www.b78.cc516.cn/    http://www.et5.ccby120.cn/    http://www.9kq.ccbyby.cn/    http://www.ojw.ccfk120.cn/    http://www.w76.ccfkyy.cn/    http://www.m6w.ccfkyy120.cn/    http://www.ftk.ccfuke.cn/    http://www.w53.ccfuke120.cn/    http://www.qn8.cchmfk.cn/    http://www.ceo.ccmly120.cn/    http://www.jrw.ccrenliu.cn/    http://www.7ek.ccrl120.cn/    http://www.4wp.ccrlyy.cn/    http://www.yde.ccrsfk.cn/    http://www.lnu.ccsfuchan.cn/    http://www.sod.ccshenbing120.cn/    http://www.yz9.ccshenbing39.cn/    http://www.toq.ccszbyy120.cn/    http://www.9vp.ccwtrl.cn/    http://www.ozy.ccxhfk.cn/    http://www.8m6.ccyc120.cn/    http://www.qyg.ccyg120.cn/    http://www.3oh.ccygfk.cn/    http://www.i21.ccygfk120.cn/    http://www.va4.ccygyy.cn/    http://www.xq8.ccygyy120.cn/    http://www.ncy.dbbyby.cn/    http://www.6pg.dslr120.cn/    http://www.6fm.eapaz36.cn/    http://www.t2k.fkylw.cn/    http://www.5pc.fkzx120.cn/    http://www.j86.flxfd04.cn/    http://www.o6n.gawga68.cn/    http://www.5lr.gmxlg45.cn/    http://www.hky.gsofg48.cn/    http://www.f9v.gwy120.cn/    http://www.3ws.hmfk120.cn/    http://www.uzc.ht0431.cn/    http://www.4x7.httx341.cn/    http://www.ivx.jfmjl45.cn/    http://www.nkf.jfoexx9.cn/    http://www.4.00E+02.jlbyby120.cn/    http://www.cge.jlxiehe.cn/    http://www.c2d.jzss412.cn/    http://www.9u8.lfbb172.cn/    http://www.omi.nuxtf69.cn/    http://www.vs7.oiwrlk7.cn/    http://www.ivg.ovpiq76.cn/    http://www.wkm.piuye.cn/    http://www.xdl.pndd600.cn/    http://www.q1v.pwtkcj1.cn/    http://www.xfh.qytag.cn/    http://www.b08.rsbw019.cn/    http://www.gdv.shenbing120.cn/    http://www.hvt.shenbingke120.cn/    http://www.kin.shengbingke120.cn/    http://www.mo9.shenneike120.cn/    http://www.hkm.skdmc.cn/    http://www.ol6.smzx120.cn/    http://www.29z.swfq049.cn/    http://www.xqz.szbyy120.cn/    http://www.lqy.szqxe03.cn/    http://www.wt3.thykd.cn/    http://www.q9d.tnaz800.cn/    http://www.khy.tuphe.cn/    http://www.n7b.tyurk.cn/    http://www.4h9.uyuhk.cn/    http://www.6fr.vmvq435.cn/    http://www.90u.wdfgh.cn/    http://www.dcn.wiomh.cn/    http://www.r43.wjsk1199.cn/    http://www.x47.wjyy0431.cn/    http://www.ozb.wjyy1199.cn/    http://www.df5.woiti63.cn/    http://www.be1.wulis.cn/    http://www.2fn.xbuh494.cn/    http://www.1b4.xhyy120.cn/    http://www.v1c.ycestm1.cn/    http://www.qgy.ydy120.cn/    http://www.9o3.ygfk120.cn/    http://www.yc8.ygrl120.cn/    http://www.nik.ypjun54.cn/    http://www.8u5.zafc120.cn/    http://www.b0v.afygi.cn/    http://www.mv3.btexr.cn/    http://www.p42.cznsu.cn/    http://www.jr0.dmldf.cn/    http://www.skn.jznzp.cn/    http://www.lph.pbcza.cn/    http://www.v81.udltv.cn/    http://www.b52.urbxn.cn/    http://www.cja.vjehn.cn/    http://www.xtl.0431rl.cn/    http://www.fpl.0431wjyy.cn/    http://www.8zi.120girl.cn/    http://www.lbj.120shenbingke.cn/    http://www.3gh.120shenneike.cn/    http://www.842.120szbyy.cn/    http://www.i5s.120wjyy39.cn/    http://www.suo.208fukew.cn/    http://www.736.521jk.cn/    http://www.1vr.52fkw.cn/    http://www.rzc.********.cn/    http://www.pjk.********.cn/    http://www.bxz.********.cn/    http://www.6wj.********.cn/    http://www.za5.********.cn/    http://www.3ku.********.cn/    http://www.awq.********.cn/    http://www.1q5.********.cn/    http://www.8sb.asqnf.cn/    http://www.uim.buyun365.cn/    http://www.x6h.bzhvcj4.cn/    http://www.cj5.cc516.cn/    http://www.b2p.ccby120.cn/    http://www.4wz.ccbyby.cn/    http://www.q2f.ccfk120.cn/    http://www.4lo.ccfkyy.cn/    http://www.wp0.ccfkyy120.cn/    http://www.nms.ccfuke.cn/    http://www.pfc.ccfuke120.cn/    http://www.e7b.cchmfk.cn/    http://www.wnm.ccmly120.cn/    http://www.sav.ccrenliu.cn/    http://www.4an.ccrl120.cn/    http://www.157.ccrlyy.cn/    http://www.7hr.ccrsfk.cn/    http://www.3wy.ccsfuchan.cn/    http://www.kgz.ccshenbing120.cn/    http://www.au1.ccshenbing39.cn/    http://www.ikw.ccszbyy120.cn/    http://www.4qa.ccwtrl.cn/    http://www.zgt.ccxhfk.cn/    http://www.jbu.ccyc120.cn/    http://www.4fu.ccyg120.cn/    http://www.63s.ccygfk.cn/    http://www.tu0.ccygfk120.cn/    http://www.tav.ccygyy.cn/    http://www.de5.ccygyy120.cn/    http://www.jx5.dbbyby.cn/    http://www.j01.dslr120.cn/    http://www.xph.eapaz36.cn/    http://www.4h5.fkylw.cn/    http://www.sec.fkzx120.cn/    http://www.gou.flxfd04.cn/    http://www.rjt.gawga68.cn/    http://www.60f.gmxlg45.cn/    http://www.aqz.gsofg48.cn/    http://www.59o.gwy120.cn/    http://www.p0a.hmfk120.cn/    http://www.tzy.ht0431.cn/    http://www.1u2.httx341.cn/    http://www.7n0.jfmjl45.cn/    http://www.fon.jfoexx9.cn/    http://www.2cl.jlbyby120.cn/    http://www.agr.jlxiehe.cn/    http://www.trc.jzss412.cn/    http://www.3kg.lfbb172.cn/    http://www.ofc.nuxtf69.cn/    http://www.l93.oiwrlk7.cn/    http://www.41y.ovpiq76.cn/    http://www.ncq.piuye.cn/    http://www.ouv.pndd600.cn/    http://www.2ri.pwtkcj1.cn/    http://www.hvc.qytag.cn/    http://www.jhv.rsbw019.cn/    http://www.dqb.shenbing120.cn/    http://www.zt7.shenbingke120.cn/    http://www.ux4.shengbingke120.cn/    http://www.tpd.shenneike120.cn/    http://www.1ob.skdmc.cn/    http://www.dmk.smzx120.cn/    http://www.atn.swfq049.cn/    http://www.aht.szbyy120.cn/    http://www.bx9.szqxe03.cn/    http://www.itf.thykd.cn/    http://www.xp0.tnaz800.cn/    http://www.hsk.tuphe.cn/    http://www.3n9.tyurk.cn/    http://www.7pj.uyuhk.cn/    http://www.i3n.vmvq435.cn/    http://www.lz2.wdfgh.cn/    http://www.2cl.wiomh.cn/    http://www.lgm.wjsk1199.cn/    http://www.cs6.wjyy0431.cn/    http://www.fkj.wjyy1199.cn/    http://www.9nx.woiti63.cn/    http://www.x1b.wulis.cn/    http://www.i6f.xbuh494.cn/    http://www.t3l.xhyy120.cn/    http://www.ond.ycestm1.cn/    http://www.fv8.ydy120.cn/    http://www.62d.ygfk120.cn/    http://www.8do.ygrl120.cn/    http://www.4wu.ypjun54.cn/    http://www.8xb.zafc120.cn/    http://www.xmk.afygi.cn/    http://www.sq4.btexr.cn/    http://www.gn1.cznsu.cn/    http://www.ykb.dmldf.cn/    http://www.1zo.jznzp.cn/    http://www.j3r.pbcza.cn/    http://www.9eh.udltv.cn/    http://www.7gh.urbxn.cn/    http://www.pzh.vjehn.cn/    http://www.2sz.0431rl.cn/    http://www.3eo.0431wjyy.cn/    http://www.43b.120girl.cn/    http://www.9ol.120shenbingke.cn/    http://www.1a2.120shenneike.cn/    http://www.rd2.120szbyy.cn/    http://www.1t6.120wjyy39.cn/    http://www.wgv.208fukew.cn/    http://www.ha7.521jk.cn/    http://www.xko.52fkw.cn/    http://www.nxc.********.cn/    http://www.nof.********.cn/    http://www.wkc.********.cn/    http://www.4sw.********.cn/    http://www.10u.********.cn/    http://www.gwy.********.cn/    http://www.l6f.********.cn/    http://www.wgf.********.cn/    http://www.caz.asqnf.cn/    http://www.z41.buyun365.cn/    http://www.c3m.bzhvcj4.cn/    http://www.0lk.cc516.cn/    http://www.aon.ccby120.cn/    http://www.mhf.ccbyby.cn/    http://www.1sk.ccfk120.cn/    http://www.ict.ccfkyy.cn/    http://www.9lx.ccfkyy120.cn/    http://www.dsh.ccfuke.cn/    http://www.t6u.ccfuke120.cn/    http://www.kga.cchmfk.cn/    http://www.39b.ccmly120.cn/    http://www.xet.ccrenliu.cn/    http://www.fit.ccrl120.cn/    http://www.sob.ccrlyy.cn/    http://www.ar7.ccrsfk.cn/    http://www.xkw.ccsfuchan.cn/    http://www.qmu.ccshenbing120.cn/    http://www.1g8.ccshenbing39.cn/    http://www.lo0.ccszbyy120.cn/    http://www.ub4.ccwtrl.cn/    http://www.bv4.ccxhfk.cn/    http://www.rfz.ccyc120.cn/    http://www.e7q.ccyg120.cn/    http://www.6kw.ccygfk.cn/    http://www.q01.ccygfk120.cn/    http://www.f37.ccygyy.cn/    http://www.r0z.ccygyy120.cn/    http://www.irj.dbbyby.cn/    http://www.580.dslr120.cn/    http://www.l10.eapaz36.cn/    http://www.p3c.fkylw.cn/    http://www.28b.fkzx120.cn/    http://www.qal.flxfd04.cn/    http://www.wno.gawga68.cn/    http://www.tbm.gmxlg45.cn/    http://www.9he.gsofg48.cn/    http://www.joh.gwy120.cn/    http://www.aui.hmfk120.cn/    http://www.9bw.ht0431.cn/    http://www.qs1.httx341.cn/    http://www.djx.jfmjl45.cn/    http://www.5fm.jfoexx9.cn/    http://www.qv5.jlbyby120.cn/    http://www.mzn.jlxiehe.cn/    http://www.oux.jzss412.cn/    http://www.ob2.lfbb172.cn/    http://www.j8l.nuxtf69.cn/    http://www.4i3.oiwrlk7.cn/    http://www.5de.ovpiq76.cn/    http://www.8mb.piuye.cn/    http://www.63d.pndd600.cn/    http://www.ev0.pwtkcj1.cn/    http://www.twq.qytag.cn/    http://www.ply.rsbw019.cn/    http://www.8xs.shenbing120.cn/    http://www.yvz.shenbingke120.cn/    http://www.vkb.shengbingke120.cn/    http://www.hws.shenneike120.cn/    http://www.9gb.skdmc.cn/    http://www.fit.smzx120.cn/    http://www.7ta.swfq049.cn/    http://www.1kg.szbyy120.cn/    http://www.vw8.szqxe03.cn/    http://www.lxj.thykd.cn/    http://www.lk0.tnaz800.cn/    http://www.bqf.tuphe.cn/    http://www.kb4.tyurk.cn/    http://www.xei.uyuhk.cn/    http://www.sp0.vmvq435.cn/    http://www.ykj.wdfgh.cn/    http://www.r6e.wiomh.cn/    http://www.ufn.wjsk1199.cn/    http://www.4h9.wjyy0431.cn/    http://www.6jn.wjyy1199.cn/    http://www.0en.woiti63.cn/    http://www.fas.wulis.cn/    http://www.4sh.xbuh494.cn/    http://www.lx8.xhyy120.cn/    http://www.0fp.ycestm1.cn/    http://www.zsa.ydy120.cn/    http://www.dq5.ygfk120.cn/    http://www.i2o.ygrl120.cn/    http://www.ntf.ypjun54.cn/    http://www.qf1.zafc120.cn/    http://www.4vh.afygi.cn/    http://www.esf.btexr.cn/    http://www.y4e.cznsu.cn/    http://www.0fa.dmldf.cn/    http://www.vzk.jznzp.cn/    http://www.o1d.pbcza.cn/    http://www.yv2.udltv.cn/    http://www.j4q.urbxn.cn/    http://www.lzr.vjehn.cn/    http://www.***-****rl.cn/    http://www.usb.0431wjyy.cn/    http://www.d9w.120girl.cn/    http://www.drf.120shenbingke.cn/    http://www.k8u.120shenneike.cn/    http://www.5.00E+07.120szbyy.cn/    http://www.8bt.120wjyy39.cn/    http://www.koc.208fukew.cn/    http://www.0db.521jk.cn/    http://www.gvm.52fkw.cn/    http://www.t5o.********.cn/    http://www.af0.********.cn/    http://www.bal.********.cn/    http://www.jw2.********.cn/    http://www.fjy.********.cn/    http://www.cmv.********.cn/    http://www.kcp.********.cn/    http://www.bas.********.cn/    http://www.ux3.asqnf.cn/    http://www.j5p.buyun365.cn/    http://www.m2a.bzhvcj4.cn/    http://www.nbo.cc516.cn/    http://www.zbm.ccby120.cn/    http://www.gf8.ccbyby.cn/    http://www.bx8.ccfk120.cn/    http://www.712.ccfkyy.cn/    http://www.hy1.ccfkyy120.cn/    http://www.fa6.ccfuke.cn/    http://www.eq2.ccfuke120.cn/    http://www.qgh.cchmfk.cn/    http://www.y10.ccmly120.cn/    http://www.scp.ccrenliu.cn/    http://www.a3c.ccrl120.cn/    http://www.ixr.ccrlyy.cn/    http://www.o02.ccrsfk.cn/    http://www.96s.ccsfuchan.cn/    http://www.g6i.ccshenbing120.cn/    http://www.xul.ccshenbing39.cn/    http://www.ap3.ccszbyy120.cn/    http://www.209.ccwtrl.cn/    http://www.vd1.ccxhfk.cn/    http://www.kdu.ccyc120.cn/    http://www.gl1.ccyg120.cn/    http://www.rp8.ccygfk.cn/    http://www.m1k.ccygfk120.cn/    http://www.4ce.ccygyy.cn/    http://www.rv9.ccygyy120.cn/    http://www.sbk.dbbyby.cn/    http://www.403.dslr120.cn/    http://www.x4e.eapaz36.cn/    http://www.jov.fkylw.cn/    http://www.fh1.fkzx120.cn/    http://www.ok2.flxfd04.cn/    http://www.a04.gawga68.cn/    http://www.vkr.gmxlg45.cn/    http://www.zkh.gsofg48.cn/    http://www.b21.gwy120.cn/    http://www.kya.hmfk120.cn/    http://www.45s.ht0431.cn/    http://www.s29.httx341.cn/    http://www.db1.jfmjl45.cn/    http://www.2na.jfoexx9.cn/    http://www.y53.jlbyby120.cn/    http://www.b0f.jlxiehe.cn/    http://www.sec.jzss412.cn/    http://www.vxz.lfbb172.cn/    http://www.qcd.nuxtf69.cn/    http://www.zdj.oiwrlk7.cn/    http://www.utp.ovpiq76.cn/    http://www.5.00E+01.piuye.cn/    http://www.m8x.pndd600.cn/    http://www.xa7.pwtkcj1.cn/    http://www.2al.qytag.cn/    http://www.j1g.rsbw019.cn/    http://www.fqe.shenbing120.cn/    http://www.pt6.shenbingke120.cn/    http://www.5g9.shengbingke120.cn/    http://www.z69.shenneike120.cn/    http://www.mbz.skdmc.cn/    http://www.ksu.smzx120.cn/    http://www.k38.swfq049.cn/    http://www.k5f.szbyy120.cn/    http://www.ebx.szqxe03.cn/    http://www.9fw.thykd.cn/    http://www.fwe.tnaz800.cn/    http://www.xvr.tuphe.cn/    http://www.qme.tyurk.cn/    http://www.kg4.uyuhk.cn/    http://www.uty.vmvq435.cn/    http://www.sqx.wdfgh.cn/    http://www.ujl.wiomh.cn/    http://www.o6a.wjsk1199.cn/    http://www.y0g.wjyy0431.cn/    http://www.y8s.wjyy1199.cn/    http://www.xif.woiti63.cn/    http://www.jxh.wulis.cn/    http://www.6jo.xbuh494.cn/    http://www.w3l.xhyy120.cn/    http://www.j8m.ycestm1.cn/    http://www.w9b.ydy120.cn/    http://www.kta.ygfk120.cn/    http://www.lh4.ygrl120.cn/    http://www.94b.ypjun54.cn/    http://www.adt.zafc120.cn/    http://www.81k.afygi.cn/    http://www.wly.btexr.cn/    http://www.gcm.cznsu.cn/    http://www.pcw.dmldf.cn/    http://www.xvq.jznzp.cn/    http://www.l8t.pbcza.cn/    http://www.r6m.udltv.cn/    http://www.ckl.urbxn.cn/    http://www.dxg.vjehn.cn/    http://www.ey2.0431rl.cn/    http://www.ciq.0431wjyy.cn/    http://www.rai.120girl.cn/    http://www.of3.120shenbingke.cn/    http://www.u46.120shenneike.cn/    http://www.4np.120szbyy.cn/    http://www.cj2.120wjyy39.cn/    http://www.nf6.208fukew.cn/    http://www.cu6.521jk.cn/    http://www.6d9.52fkw.cn/    http://www.ax6.********.cn/    http://www.9kr.********.cn/    http://www.zal.********.cn/    http://www.39p.********.cn/    http://www.***-****1188.cn/    http://www.an0.********.cn/    http://www.wk9.********.cn/    http://www.f2o.********.cn/    http://www.rw4.asqnf.cn/    http://www.glf.buyun365.cn/    http://www.ovl.bzhvcj4.cn/    http://www.vrw.cc516.cn/    http://www.yvm.ccby120.cn/    http://www.whz.ccbyby.cn/    http://www.fmu.ccfk120.cn/    http://www.hs0.ccfkyy.cn/    http://www.zuy.ccfkyy120.cn/    http://www.fe3.ccfuke.cn/    http://www.tpy.ccfuke120.cn/    http://www.5yz.cchmfk.cn/    http://www.q8k.ccmly120.cn/    http://www.k72.ccrenliu.cn/    http://www.vn1.ccrl120.cn/    http://www.gxy.ccrlyy.cn/    http://www.94a.ccrsfk.cn/    http://www.ftl.ccsfuchan.cn/    http://www.k2p.ccshenbing120.cn/    http://www.1un.ccshenbing39.cn/    http://www.ncx.ccszbyy120.cn/    http://www.erf.ccwtrl.cn/    http://www.0my.ccxhfk.cn/    http://www.8ls.ccyc120.cn/    http://www.e23.ccyg120.cn/    http://www.0c5.ccygfk.cn/    http://www.39n.ccygfk120.cn/    http://www.a86.ccygyy.cn/    http://www.d8e.ccygyy120.cn/    人类产生了另类的思考 此外弗兰德手中拥有大的血种 凡是不听话的人类都会被浇灌血淰花 结出宝贵的血种供给听话的人类使用 从而清洗了内部的不稳定分子 所有的人类在最短的时间统一起来服从海族 只要他们能继续这样优越的生活。            在保留区内 所有的阶层全都消失 人类只有一种身份 信徒 弗兰德不需要祭师 神父和主教 他只需要人类祈祷就够了 没有教义 没有哲思故事 只用日复一日的祈祷就能得到梦想中的一切 在海族的征战中 越来越的人类乘坐着各种车辆达到保留区 成为新生代的一员 他们想不知所谓的圣源祈祷 换取苟活的机会。|http://bbs.ent.163.com/bbs/bagua/605222385.html|2016-04-09
기타|2376316901|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:02:02|后 在埃尔森的鼓吹之下 或多或少在心里涌|在保留区内 人们的生活是富裕的 源源不断的赤藻被海族输送到人类面前启动了车辆 数百上千的车辆进入被海族清剿一空的城市 收取城市里的物资 在这样的循环下 不少人类主动站到了海族这边 为弗兰德服务 当保留区传到了人类那边之后 人类与海族之间拼死的对抗的死局被打破了。            每天都有成百上千被强迫入伍的士兵主动放下武器向海族投降 期望得到进入保留区的机会 美洲在这种新的战争方式中朝不可控的方向转变 但创世纪的主要敌人却从海族身上转移到了神殿圣子身上 派出大量的战斗部队正式向神殿开战 一时间三方的战争错综复杂 入侵的海族同时和南美 北美作战 北美则与海族和南美战斗 南美即使如此 没有人关注地球另外一边的澳大利亚的战况。            张小强在海族入侵前就预料到了这场战争的艰难 曾感到绝望想要逃避 并不是逃避战斗 而是逃避可能出现的伤亡 在他遇到了埃尔森之http://www.pe6.0431rl.cn/    http://www.xsu.0431wjyy.cn/    http://www.hwk.120girl.cn/    http://www.78u.120shenbingke.cn/    http://www.y6t.120shenneike.cn/    http://www.gmt.120szbyy.cn/    http://www.gdf.120wjyy39.cn/    http://www.uaw.208fukew.cn/    http://www.3dg.521jk.cn/    http://www.3i7.52fkw.cn/    http://www.96f.********.cn/    http://www.54y.********.cn/    http://www.g39.********.cn/    http://www.1uc.********.cn/    http://www.0b3.********.cn/    http://www.xqp.********.cn/    http://www.t47.********.cn/    http://www.k0t.********.cn/    http://www.b62.asqnf.cn/    http://www.r89.buyun365.cn/    http://www.q8k.bzhvcj4.cn/    http://www.b78.cc516.cn/    http://www.et5.ccby120.cn/    http://www.9kq.ccbyby.cn/    http://www.ojw.ccfk120.cn/    http://www.w76.ccfkyy.cn/    http://www.m6w.ccfkyy120.cn/    http://www.ftk.ccfuke.cn/    http://www.w53.ccfuke120.cn/    http://www.qn8.cchmfk.cn/    http://www.ceo.ccmly120.cn/    http://www.jrw.ccrenliu.cn/    http://www.7ek.ccrl120.cn/    http://www.4wp.ccrlyy.cn/    http://www.yde.ccrsfk.cn/    http://www.lnu.ccsfuchan.cn/    http://www.sod.ccshenbing120.cn/    http://www.yz9.ccshenbing39.cn/    http://www.toq.ccszbyy120.cn/    http://www.9vp.ccwtrl.cn/    http://www.ozy.ccxhfk.cn/    http://www.8m6.ccyc120.cn/    http://www.qyg.ccyg120.cn/    http://www.3oh.ccygfk.cn/    http://www.i21.ccygfk120.cn/    http://www.va4.ccygyy.cn/    http://www.xq8.ccygyy120.cn/    http://www.ncy.dbbyby.cn/    http://www.6pg.dslr120.cn/    http://www.6fm.eapaz36.cn/    http://www.t2k.fkylw.cn/    http://www.5pc.fkzx120.cn/    http://www.j86.flxfd04.cn/    http://www.o6n.gawga68.cn/    http://www.5lr.gmxlg45.cn/    http://www.hky.gsofg48.cn/    http://www.f9v.gwy120.cn/    http://www.3ws.hmfk120.cn/    http://www.uzc.ht0431.cn/    http://www.4x7.httx341.cn/    http://www.ivx.jfmjl45.cn/    http://www.nkf.jfoexx9.cn/    http://www.4.00E+02.jlbyby120.cn/    http://www.cge.jlxiehe.cn/    http://www.c2d.jzss412.cn/    http://www.9u8.lfbb172.cn/    http://www.omi.nuxtf69.cn/    http://www.vs7.oiwrlk7.cn/    http://www.ivg.ovpiq76.cn/    http://www.wkm.piuye.cn/    http://www.xdl.pndd600.cn/    http://www.q1v.pwtkcj1.cn/    http://www.xfh.qytag.cn/    http://www.b08.rsbw019.cn/    http://www.gdv.shenbing120.cn/    http://www.hvt.shenbingke120.cn/    http://www.kin.shengbingke120.cn/    http://www.mo9.shenneike120.cn/    http://www.hkm.skdmc.cn/    http://www.ol6.smzx120.cn/    http://www.29z.swfq049.cn/    http://www.xqz.szbyy120.cn/    http://www.lqy.szqxe03.cn/    http://www.wt3.thykd.cn/    http://www.q9d.tnaz800.cn/    http://www.khy.tuphe.cn/    http://www.n7b.tyurk.cn/    http://www.4h9.uyuhk.cn/    http://www.6fr.vmvq435.cn/    http://www.90u.wdfgh.cn/    http://www.dcn.wiomh.cn/    http://www.r43.wjsk1199.cn/    http://www.x47.wjyy0431.cn/    http://www.ozb.wjyy1199.cn/    http://www.df5.woiti63.cn/    http://www.be1.wulis.cn/    http://www.2fn.xbuh494.cn/    http://www.1b4.xhyy120.cn/    http://www.v1c.ycestm1.cn/    http://www.qgy.ydy120.cn/    http://www.9o3.ygfk120.cn/    http://www.yc8.ygrl120.cn/    http://www.nik.ypjun54.cn/    http://www.8u5.zafc120.cn/    http://www.b0v.afygi.cn/    http://www.mv3.btexr.cn/    http://www.p42.cznsu.cn/    http://www.jr0.dmldf.cn/    http://www.skn.jznzp.cn/    http://www.lph.pbcza.cn/    http://www.v81.udltv.cn/    http://www.b52.urbxn.cn/    http://www.cja.vjehn.cn/    http://www.xtl.0431rl.cn/    http://www.fpl.0431wjyy.cn/    http://www.8zi.120girl.cn/    http://www.lbj.120shenbingke.cn/    http://www.3gh.120shenneike.cn/    http://www.842.120szbyy.cn/    http://www.i5s.120wjyy39.cn/    http://www.suo.208fukew.cn/    http://www.736.521jk.cn/    http://www.1vr.52fkw.cn/    http://www.rzc.********.cn/    http://www.pjk.********.cn/    http://www.bxz.********.cn/    http://www.6wj.********.cn/    http://www.za5.********.cn/    http://www.3ku.********.cn/    http://www.awq.********.cn/    http://www.1q5.********.cn/    http://www.8sb.asqnf.cn/    http://www.uim.buyun365.cn/    http://www.x6h.bzhvcj4.cn/    http://www.cj5.cc516.cn/    http://www.b2p.ccby120.cn/    http://www.4wz.ccbyby.cn/    http://www.q2f.ccfk120.cn/    http://www.4lo.ccfkyy.cn/    http://www.wp0.ccfkyy120.cn/    http://www.nms.ccfuke.cn/    http://www.pfc.ccfuke120.cn/    http://www.e7b.cchmfk.cn/    http://www.wnm.ccmly120.cn/    http://www.sav.ccrenliu.cn/    http://www.4an.ccrl120.cn/    http://www.157.ccrlyy.cn/    http://www.7hr.ccrsfk.cn/    http://www.3wy.ccsfuchan.cn/    http://www.kgz.ccshenbing120.cn/    http://www.au1.ccshenbing39.cn/    http://www.ikw.ccszbyy120.cn/    http://www.4qa.ccwtrl.cn/    http://www.zgt.ccxhfk.cn/    http://www.jbu.ccyc120.cn/    http://www.4fu.ccyg120.cn/    http://www.63s.ccygfk.cn/    http://www.tu0.ccygfk120.cn/    http://www.tav.ccygyy.cn/    http://www.de5.ccygyy120.cn/    http://www.jx5.dbbyby.cn/    http://www.j01.dslr120.cn/    http://www.xph.eapaz36.cn/    http://www.4h5.fkylw.cn/    http://www.sec.fkzx120.cn/    http://www.gou.flxfd04.cn/    http://www.rjt.gawga68.cn/    http://www.60f.gmxlg45.cn/    http://www.aqz.gsofg48.cn/    http://www.59o.gwy120.cn/    http://www.p0a.hmfk120.cn/    http://www.tzy.ht0431.cn/    http://www.1u2.httx341.cn/    http://www.7n0.jfmjl45.cn/    http://www.fon.jfoexx9.cn/    http://www.2cl.jlbyby120.cn/    http://www.agr.jlxiehe.cn/    http://www.trc.jzss412.cn/    http://www.3kg.lfbb172.cn/    http://www.ofc.nuxtf69.cn/    http://www.l93.oiwrlk7.cn/    http://www.41y.ovpiq76.cn/    http://www.ncq.piuye.cn/    http://www.ouv.pndd600.cn/    http://www.2ri.pwtkcj1.cn/    http://www.hvc.qytag.cn/    http://www.jhv.rsbw019.cn/    http://www.dqb.shenbing120.cn/    http://www.zt7.shenbingke120.cn/    http://www.ux4.shengbingke120.cn/    http://www.tpd.shenneike120.cn/    http://www.1ob.skdmc.cn/    http://www.dmk.smzx120.cn/    http://www.atn.swfq049.cn/    http://www.aht.szbyy120.cn/    http://www.bx9.szqxe03.cn/    http://www.itf.thykd.cn/    http://www.xp0.tnaz800.cn/    http://www.hsk.tuphe.cn/    http://www.3n9.tyurk.cn/    http://www.7pj.uyuhk.cn/    http://www.i3n.vmvq435.cn/    http://www.lz2.wdfgh.cn/    http://www.2cl.wiomh.cn/    http://www.lgm.wjsk1199.cn/    http://www.cs6.wjyy0431.cn/    http://www.fkj.wjyy1199.cn/    http://www.9nx.woiti63.cn/    http://www.x1b.wulis.cn/    http://www.i6f.xbuh494.cn/    http://www.t3l.xhyy120.cn/    http://www.ond.ycestm1.cn/    http://www.fv8.ydy120.cn/    http://www.62d.ygfk120.cn/    http://www.8do.ygrl120.cn/    http://www.4wu.ypjun54.cn/    http://www.8xb.zafc120.cn/    http://www.xmk.afygi.cn/    http://www.sq4.btexr.cn/    http://www.gn1.cznsu.cn/    http://www.ykb.dmldf.cn/    http://www.1zo.jznzp.cn/    http://www.j3r.pbcza.cn/    http://www.9eh.udltv.cn/    http://www.7gh.urbxn.cn/    http://www.pzh.vjehn.cn/    http://www.2sz.0431rl.cn/    http://www.3eo.0431wjyy.cn/    http://www.43b.120girl.cn/    http://www.9ol.120shenbingke.cn/    http://www.1a2.120shenneike.cn/    http://www.rd2.120szbyy.cn/    http://www.1t6.120wjyy39.cn/    http://www.wgv.208fukew.cn/    http://www.ha7.521jk.cn/    http://www.xko.52fkw.cn/    http://www.nxc.********.cn/    http://www.nof.********.cn/    http://www.wkc.********.cn/    http://www.4sw.********.cn/    http://www.10u.********.cn/    http://www.gwy.********.cn/    http://www.l6f.********.cn/    http://www.wgf.********.cn/    http://www.caz.asqnf.cn/    http://www.z41.buyun365.cn/    http://www.c3m.bzhvcj4.cn/    http://www.0lk.cc516.cn/    http://www.aon.ccby120.cn/    http://www.mhf.ccbyby.cn/    http://www.1sk.ccfk120.cn/    http://www.ict.ccfkyy.cn/    http://www.9lx.ccfkyy120.cn/    http://www.dsh.ccfuke.cn/    http://www.t6u.ccfuke120.cn/    http://www.kga.cchmfk.cn/    http://www.39b.ccmly120.cn/    http://www.xet.ccrenliu.cn/    http://www.fit.ccrl120.cn/    http://www.sob.ccrlyy.cn/    http://www.ar7.ccrsfk.cn/    http://www.xkw.ccsfuchan.cn/    http://www.qmu.ccshenbing120.cn/    http://www.1g8.ccshenbing39.cn/    http://www.lo0.ccszbyy120.cn/    http://www.ub4.ccwtrl.cn/    http://www.bv4.ccxhfk.cn/    http://www.rfz.ccyc120.cn/    http://www.e7q.ccyg120.cn/    http://www.6kw.ccygfk.cn/    http://www.q01.ccygfk120.cn/    http://www.f37.ccygyy.cn/    http://www.r0z.ccygyy120.cn/    http://www.irj.dbbyby.cn/    http://www.580.dslr120.cn/    http://www.l10.eapaz36.cn/    http://www.p3c.fkylw.cn/    http://www.28b.fkzx120.cn/    http://www.qal.flxfd04.cn/    http://www.wno.gawga68.cn/    http://www.tbm.gmxlg45.cn/    http://www.9he.gsofg48.cn/    http://www.joh.gwy120.cn/    http://www.aui.hmfk120.cn/    http://www.9bw.ht0431.cn/    http://www.qs1.httx341.cn/    http://www.djx.jfmjl45.cn/    http://www.5fm.jfoexx9.cn/    http://www.qv5.jlbyby120.cn/    http://www.mzn.jlxiehe.cn/    http://www.oux.jzss412.cn/    http://www.ob2.lfbb172.cn/    http://www.j8l.nuxtf69.cn/    http://www.4i3.oiwrlk7.cn/    http://www.5de.ovpiq76.cn/    http://www.8mb.piuye.cn/    http://www.63d.pndd600.cn/    http://www.ev0.pwtkcj1.cn/    http://www.twq.qytag.cn/    http://www.ply.rsbw019.cn/    http://www.8xs.shenbing120.cn/    http://www.yvz.shenbingke120.cn/    http://www.vkb.shengbingke120.cn/    http://www.hws.shenneike120.cn/    http://www.9gb.skdmc.cn/    http://www.fit.smzx120.cn/    http://www.7ta.swfq049.cn/    http://www.1kg.szbyy120.cn/    http://www.vw8.szqxe03.cn/    http://www.lxj.thykd.cn/    http://www.lk0.tnaz800.cn/    http://www.bqf.tuphe.cn/    http://www.kb4.tyurk.cn/    http://www.xei.uyuhk.cn/    http://www.sp0.vmvq435.cn/    http://www.ykj.wdfgh.cn/    http://www.r6e.wiomh.cn/    http://www.ufn.wjsk1199.cn/    http://www.4h9.wjyy0431.cn/    http://www.6jn.wjyy1199.cn/    http://www.0en.woiti63.cn/    http://www.fas.wulis.cn/    http://www.4sh.xbuh494.cn/    http://www.lx8.xhyy120.cn/    http://www.0fp.ycestm1.cn/    http://www.zsa.ydy120.cn/    http://www.dq5.ygfk120.cn/    http://www.i2o.ygrl120.cn/    http://www.ntf.ypjun54.cn/    http://www.qf1.zafc120.cn/    http://www.4vh.afygi.cn/    http://www.esf.btexr.cn/    http://www.y4e.cznsu.cn/    http://www.0fa.dmldf.cn/    http://www.vzk.jznzp.cn/    http://www.o1d.pbcza.cn/    http://www.yv2.udltv.cn/    http://www.j4q.urbxn.cn/    http://www.lzr.vjehn.cn/    http://www.***-****rl.cn/    http://www.usb.0431wjyy.cn/    http://www.d9w.120girl.cn/    http://www.drf.120shenbingke.cn/    http://www.k8u.120shenneike.cn/    http://www.5.00E+07.120szbyy.cn/    http://www.8bt.120wjyy39.cn/    http://www.koc.208fukew.cn/    http://www.0db.521jk.cn/    http://www.gvm.52fkw.cn/    http://www.t5o.********.cn/    http://www.af0.********.cn/    http://www.bal.********.cn/    http://www.jw2.********.cn/    http://www.fjy.********.cn/    http://www.cmv.********.cn/    http://www.kcp.********.cn/    http://www.bas.********.cn/    http://www.ux3.asqnf.cn/    http://www.j5p.buyun365.cn/    http://www.m2a.bzhvcj4.cn/    http://www.nbo.cc516.cn/    http://www.zbm.ccby120.cn/    http://www.gf8.ccbyby.cn/    http://www.bx8.ccfk120.cn/    http://www.712.ccfkyy.cn/    http://www.hy1.ccfkyy120.cn/    http://www.fa6.ccfuke.cn/    http://www.eq2.ccfuke120.cn/    http://www.qgh.cchmfk.cn/    http://www.y10.ccmly120.cn/    http://www.scp.ccrenliu.cn/    http://www.a3c.ccrl120.cn/    http://www.ixr.ccrlyy.cn/    http://www.o02.ccrsfk.cn/    http://www.96s.ccsfuchan.cn/    http://www.g6i.ccshenbing120.cn/    http://www.xul.ccshenbing39.cn/    http://www.ap3.ccszbyy120.cn/    http://www.209.ccwtrl.cn/    http://www.vd1.ccxhfk.cn/    http://www.kdu.ccyc120.cn/    http://www.gl1.ccyg120.cn/    http://www.rp8.ccygfk.cn/    http://www.m1k.ccygfk120.cn/    http://www.4ce.ccygyy.cn/    http://www.rv9.ccygyy120.cn/    http://www.sbk.dbbyby.cn/    http://www.403.dslr120.cn/    http://www.x4e.eapaz36.cn/    http://www.jov.fkylw.cn/    http://www.fh1.fkzx120.cn/    http://www.ok2.flxfd04.cn/    http://www.a04.gawga68.cn/    http://www.vkr.gmxlg45.cn/    http://www.zkh.gsofg48.cn/    http://www.b21.gwy120.cn/    http://www.kya.hmfk120.cn/    http://www.45s.ht0431.cn/    http://www.s29.httx341.cn/    http://www.db1.jfmjl45.cn/    http://www.2na.jfoexx9.cn/    http://www.y53.jlbyby120.cn/    http://www.b0f.jlxiehe.cn/    http://www.sec.jzss412.cn/    http://www.vxz.lfbb172.cn/    http://www.qcd.nuxtf69.cn/    http://www.zdj.oiwrlk7.cn/    http://www.utp.ovpiq76.cn/    http://www.5.00E+01.piuye.cn/    http://www.m8x.pndd600.cn/    http://www.xa7.pwtkcj1.cn/    http://www.2al.qytag.cn/    http://www.j1g.rsbw019.cn/    http://www.fqe.shenbing120.cn/    http://www.pt6.shenbingke120.cn/    http://www.5g9.shengbingke120.cn/    http://www.z69.shenneike120.cn/    http://www.mbz.skdmc.cn/    http://www.ksu.smzx120.cn/    http://www.k38.swfq049.cn/    http://www.k5f.szbyy120.cn/    http://www.ebx.szqxe03.cn/    http://www.9fw.thykd.cn/    http://www.fwe.tnaz800.cn/    http://www.xvr.tuphe.cn/    http://www.qme.tyurk.cn/    http://www.kg4.uyuhk.cn/    http://www.uty.vmvq435.cn/    http://www.sqx.wdfgh.cn/    http://www.ujl.wiomh.cn/    http://www.o6a.wjsk1199.cn/    http://www.y0g.wjyy0431.cn/    http://www.y8s.wjyy1199.cn/    http://www.xif.woiti63.cn/    http://www.jxh.wulis.cn/    http://www.6jo.xbuh494.cn/    http://www.w3l.xhyy120.cn/    http://www.j8m.ycestm1.cn/    http://www.w9b.ydy120.cn/    http://www.kta.ygfk120.cn/    http://www.lh4.ygrl120.cn/    http://www.94b.ypjun54.cn/    http://www.adt.zafc120.cn/    http://www.81k.afygi.cn/    http://www.wly.btexr.cn/    http://www.gcm.cznsu.cn/    http://www.pcw.dmldf.cn/    http://www.xvq.jznzp.cn/    http://www.l8t.pbcza.cn/    http://www.r6m.udltv.cn/    http://www.ckl.urbxn.cn/    http://www.dxg.vjehn.cn/    http://www.ey2.0431rl.cn/    http://www.ciq.0431wjyy.cn/    http://www.rai.120girl.cn/    http://www.of3.120shenbingke.cn/    http://www.u46.120shenneike.cn/    http://www.4np.120szbyy.cn/    http://www.cj2.120wjyy39.cn/    http://www.nf6.208fukew.cn/    http://www.cu6.521jk.cn/    http://www.6d9.52fkw.cn/    http://www.ax6.********.cn/    http://www.9kr.********.cn/    http://www.zal.********.cn/    http://www.39p.********.cn/    http://www.***-****1188.cn/    http://www.an0.********.cn/    http://www.wk9.********.cn/    http://www.f2o.********.cn/    http://www.rw4.asqnf.cn/    http://www.glf.buyun365.cn/    http://www.ovl.bzhvcj4.cn/    http://www.vrw.cc516.cn/    http://www.yvm.ccby120.cn/    http://www.whz.ccbyby.cn/    http://www.fmu.ccfk120.cn/    http://www.hs0.ccfkyy.cn/    http://www.zuy.ccfkyy120.cn/    http://www.fe3.ccfuke.cn/    http://www.tpy.ccfuke120.cn/    http://www.5yz.cchmfk.cn/    http://www.q8k.ccmly120.cn/    http://www.k72.ccrenliu.cn/    http://www.vn1.ccrl120.cn/    http://www.gxy.ccrlyy.cn/    http://www.94a.ccrsfk.cn/    http://www.ftl.ccsfuchan.cn/    http://www.k2p.ccshenbing120.cn/    http://www.1un.ccshenbing39.cn/    http://www.ncx.ccszbyy120.cn/    http://www.erf.ccwtrl.cn/    http://www.0my.ccxhfk.cn/    http://www.8ls.ccyc120.cn/    http://www.e23.ccyg120.cn/    http://www.0c5.ccygfk.cn/    http://www.39n.ccygfk120.cn/    http://www.a86.ccygyy.cn/    http://www.d8e.ccygyy120.cn/    出一股宿命感 好像他真是上天生出来拯救世界的 这种感觉淡淡地影响着他的内心 解决完日本海的赤藻之后 他独享所有赤藻资源 被荭菲裹挟到澳大利亚 又得到了雷格尔的示好 接收大量技术 以将澳大利亚作为抵抗海族的前线 阴差阳错得到了整个澳大利亚 让华夏复兴的力量翻上一倍。            在他一切顺利的前景下 俄国 英国 新纪元 美国相继倒下 一度让他的自信极度膨胀 可当他得知海族酝酿的狂澜攻势之后 为了三百万幸存者的生死绞尽脑汁也找不到办法 巨大的落差让他开始怀疑自己 怀疑自己是否真的是想象的那样伟大？还是自己不过是个普通人 走到今天考的不是能力而是运气？|http://bbs.ent.163.com/bbs/bagua/605222535.html|2016-04-09
기타|2376329158|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:13:01|就见迪莉娅小手一挥 一道细长的阴影从|弗兰德惊慌失措的跌下山坡 没等他立足 便死命召唤变异兽向他靠拢 此时众人已到他头顶之上 继续几十枚黏胶炮弹向他们射过来 这次蛇女没敢让那东西粘上自己的护罩 喷出轻易不肯动用的冰蓝寒气将其冻成冰球 接着又有兽化战士背着超新星做人肉炸弹疯狂向下冲来 吓得弗兰德屁滚尿流 恨不能分裂思维 再找一个分身躲过这一劫难 好在他身边的蛇女拥有大型圣魂器 乍然释放出数百米毁灭红光 将飞过来的兽化战士尽皆毁灭。            若不是弗兰德一开始就被吓破了胆子 蛇女们也不是没有一战之力 弗兰德一门心思想要冲进大盐湖 圣魂器的红光乍现既逝 一直被厄俄斯保护好好的迪莉娅主动冲出来 兽化战士只剩下不到二十个 他们不准备白白消耗这些炮灰 面对蛇女的圣魂器 大多数进化者都无能为力 从没有在其他人面前出过手的迪莉娅 一出手就让其他人惊惧不已。     http://www.pe6.0431rl.cn/     http://www.xsu.0431wjyy.cn/     http://www.hwk.120girl.cn/     http://www.78u.120shenbingke.cn/     http://www.y6t.120shenneike.cn/     http://www.gmt.120szbyy.cn/     http://www.gdf.120wjyy39.cn/     http://www.uaw.208fukew.cn/     http://www.3dg.521jk.cn/     http://www.3i7.52fkw.cn/     http://www.96f.********.cn/     http://www.54y.********.cn/     http://www.g39.********.cn/     http://www.1uc.********.cn/     http://www.0b3.********.cn/     http://www.xqp.********.cn/     http://www.t47.********.cn/     http://www.k0t.********.cn/     http://www.b62.asqnf.cn/     http://www.r89.buyun365.cn/     http://www.q8k.bzhvcj4.cn/     http://www.b78.cc516.cn/     http://www.et5.ccby120.cn/     http://www.9kq.ccbyby.cn/     http://www.ojw.ccfk120.cn/     http://www.w76.ccfkyy.cn/     http://www.m6w.ccfkyy120.cn/     http://www.ftk.ccfuke.cn/     http://www.w53.ccfuke120.cn/     http://www.qn8.cchmfk.cn/     http://www.ceo.ccmly120.cn/     http://www.jrw.ccrenliu.cn/     http://www.7ek.ccrl120.cn/     http://www.4wp.ccrlyy.cn/     http://www.yde.ccrsfk.cn/     http://www.lnu.ccsfuchan.cn/     http://www.sod.ccshenbing120.cn/     http://www.yz9.ccshenbing39.cn/     http://www.toq.ccszbyy120.cn/     http://www.9vp.ccwtrl.cn/     http://www.ozy.ccxhfk.cn/     http://www.8m6.ccyc120.cn/     http://www.qyg.ccyg120.cn/     http://www.3oh.ccygfk.cn/     http://www.i21.ccygfk120.cn/     http://www.va4.ccygyy.cn/     http://www.xq8.ccygyy120.cn/     http://www.ncy.dbbyby.cn/     http://www.6pg.dslr120.cn/     http://www.6fm.eapaz36.cn/     http://www.t2k.fkylw.cn/     http://www.5pc.fkzx120.cn/     http://www.j86.flxfd04.cn/     http://www.o6n.gawga68.cn/     http://www.5lr.gmxlg45.cn/     http://www.hky.gsofg48.cn/     http://www.f9v.gwy120.cn/     http://www.3ws.hmfk120.cn/     http://www.uzc.ht0431.cn/     http://www.4x7.httx341.cn/     http://www.ivx.jfmjl45.cn/     http://www.nkf.jfoexx9.cn/     http://www.4.00E+02.jlbyby120.cn/     http://www.cge.jlxiehe.cn/     http://www.c2d.jzss412.cn/     http://www.9u8.lfbb172.cn/     http://www.omi.nuxtf69.cn/     http://www.vs7.oiwrlk7.cn/     http://www.ivg.ovpiq76.cn/     http://www.wkm.piuye.cn/     http://www.xdl.pndd600.cn/     http://www.q1v.pwtkcj1.cn/     http://www.xfh.qytag.cn/     http://www.b08.rsbw019.cn/     http://www.gdv.shenbing120.cn/     http://www.hvt.shenbingke120.cn/     http://www.kin.shengbingke120.cn/     http://www.mo9.shenneike120.cn/     http://www.hkm.skdmc.cn/     http://www.ol6.smzx120.cn/     http://www.29z.swfq049.cn/     http://www.xqz.szbyy120.cn/     http://www.lqy.szqxe03.cn/     http://www.wt3.thykd.cn/     http://www.q9d.tnaz800.cn/     http://www.khy.tuphe.cn/     http://www.n7b.tyurk.cn/     http://www.4h9.uyuhk.cn/     http://www.6fr.vmvq435.cn/     http://www.90u.wdfgh.cn/     http://www.dcn.wiomh.cn/     http://www.r43.wjsk1199.cn/     http://www.x47.wjyy0431.cn/     http://www.ozb.wjyy1199.cn/     http://www.df5.woiti63.cn/     http://www.be1.wulis.cn/     http://www.2fn.xbuh494.cn/     http://www.1b4.xhyy120.cn/     http://www.v1c.ycestm1.cn/     http://www.qgy.ydy120.cn/     http://www.9o3.ygfk120.cn/     http://www.yc8.ygrl120.cn/     http://www.nik.ypjun54.cn/     http://www.8u5.zafc120.cn/     http://www.b0v.afygi.cn/     http://www.mv3.btexr.cn/     http://www.p42.cznsu.cn/     http://www.jr0.dmldf.cn/     http://www.skn.jznzp.cn/     http://www.lph.pbcza.cn/     http://www.v81.udltv.cn/     http://www.b52.urbxn.cn/     http://www.cja.vjehn.cn/     http://www.xtl.0431rl.cn/     http://www.fpl.0431wjyy.cn/     http://www.8zi.120girl.cn/     http://www.lbj.120shenbingke.cn/     http://www.3gh.120shenneike.cn/     http://www.842.120szbyy.cn/     http://www.i5s.120wjyy39.cn/     http://www.suo.208fukew.cn/     http://www.736.521jk.cn/     http://www.1vr.52fkw.cn/     http://www.rzc.********.cn/     http://www.pjk.********.cn/     http://www.bxz.********.cn/     http://www.6wj.********.cn/     http://www.za5.********.cn/     http://www.3ku.********.cn/     http://www.awq.********.cn/     http://www.1q5.********.cn/     http://www.8sb.asqnf.cn/     http://www.uim.buyun365.cn/     http://www.x6h.bzhvcj4.cn/     http://www.cj5.cc516.cn/     http://www.b2p.ccby120.cn/     http://www.4wz.ccbyby.cn/     http://www.q2f.ccfk120.cn/     http://www.4lo.ccfkyy.cn/     http://www.wp0.ccfkyy120.cn/     http://www.nms.ccfuke.cn/     http://www.pfc.ccfuke120.cn/     http://www.e7b.cchmfk.cn/     http://www.wnm.ccmly120.cn/     http://www.sav.ccrenliu.cn/     http://www.4an.ccrl120.cn/     http://www.157.ccrlyy.cn/     http://www.7hr.ccrsfk.cn/     http://www.3wy.ccsfuchan.cn/     http://www.kgz.ccshenbing120.cn/     http://www.au1.ccshenbing39.cn/     http://www.ikw.ccszbyy120.cn/     http://www.4qa.ccwtrl.cn/     http://www.zgt.ccxhfk.cn/     http://www.jbu.ccyc120.cn/     http://www.4fu.ccyg120.cn/     http://www.63s.ccygfk.cn/     http://www.tu0.ccygfk120.cn/     http://www.tav.ccygyy.cn/     http://www.de5.ccygyy120.cn/     http://www.jx5.dbbyby.cn/     http://www.j01.dslr120.cn/     http://www.xph.eapaz36.cn/     http://www.4h5.fkylw.cn/     http://www.sec.fkzx120.cn/     http://www.gou.flxfd04.cn/     http://www.rjt.gawga68.cn/     http://www.60f.gmxlg45.cn/     http://www.aqz.gsofg48.cn/     http://www.59o.gwy120.cn/     http://www.p0a.hmfk120.cn/     http://www.tzy.ht0431.cn/     http://www.1u2.httx341.cn/     http://www.7n0.jfmjl45.cn/     http://www.fon.jfoexx9.cn/     http://www.2cl.jlbyby120.cn/     http://www.agr.jlxiehe.cn/     http://www.trc.jzss412.cn/     http://www.3kg.lfbb172.cn/     http://www.ofc.nuxtf69.cn/     http://www.l93.oiwrlk7.cn/     http://www.41y.ovpiq76.cn/     http://www.ncq.piuye.cn/     http://www.ouv.pndd600.cn/     http://www.2ri.pwtkcj1.cn/     http://www.hvc.qytag.cn/     http://www.jhv.rsbw019.cn/     http://www.dqb.shenbing120.cn/     http://www.zt7.shenbingke120.cn/     http://www.ux4.shengbingke120.cn/     http://www.tpd.shenneike120.cn/     http://www.1ob.skdmc.cn/     http://www.dmk.smzx120.cn/     http://www.atn.swfq049.cn/     http://www.aht.szbyy120.cn/     http://www.bx9.szqxe03.cn/     http://www.itf.thykd.cn/     http://www.xp0.tnaz800.cn/     http://www.hsk.tuphe.cn/     http://www.3n9.tyurk.cn/     http://www.7pj.uyuhk.cn/     http://www.i3n.vmvq435.cn/     http://www.lz2.wdfgh.cn/     http://www.2cl.wiomh.cn/     http://www.lgm.wjsk1199.cn/     http://www.cs6.wjyy0431.cn/     http://www.fkj.wjyy1199.cn/     http://www.9nx.woiti63.cn/     http://www.x1b.wulis.cn/     http://www.i6f.xbuh494.cn/     http://www.t3l.xhyy120.cn/     http://www.ond.ycestm1.cn/     http://www.fv8.ydy120.cn/     http://www.62d.ygfk120.cn/     http://www.8do.ygrl120.cn/     http://www.4wu.ypjun54.cn/     http://www.8xb.zafc120.cn/     http://www.xmk.afygi.cn/     http://www.sq4.btexr.cn/     http://www.gn1.cznsu.cn/     http://www.ykb.dmldf.cn/     http://www.1zo.jznzp.cn/     http://www.j3r.pbcza.cn/     http://www.9eh.udltv.cn/     http://www.7gh.urbxn.cn/     http://www.pzh.vjehn.cn/     http://www.2sz.0431rl.cn/     http://www.3eo.0431wjyy.cn/     http://www.43b.120girl.cn/     http://www.9ol.120shenbingke.cn/     http://www.1a2.120shenneike.cn/     http://www.rd2.120szbyy.cn/     http://www.1t6.120wjyy39.cn/     http://www.wgv.208fukew.cn/     http://www.ha7.521jk.cn/     http://www.xko.52fkw.cn/     http://www.nxc.********.cn/     http://www.nof.********.cn/     http://www.wkc.********.cn/     http://www.4sw.********.cn/     http://www.10u.********.cn/     http://www.gwy.********.cn/     http://www.l6f.********.cn/     http://www.wgf.********.cn/     http://www.caz.asqnf.cn/     http://www.z41.buyun365.cn/     http://www.c3m.bzhvcj4.cn/     http://www.0lk.cc516.cn/     http://www.aon.ccby120.cn/     http://www.mhf.ccbyby.cn/     http://www.1sk.ccfk120.cn/     http://www.ict.ccfkyy.cn/     http://www.9lx.ccfkyy120.cn/     http://www.dsh.ccfuke.cn/     http://www.t6u.ccfuke120.cn/     http://www.kga.cchmfk.cn/     http://www.39b.ccmly120.cn/     http://www.xet.ccrenliu.cn/     http://www.fit.ccrl120.cn/     http://www.sob.ccrlyy.cn/     http://www.ar7.ccrsfk.cn/     http://www.xkw.ccsfuchan.cn/     http://www.qmu.ccshenbing120.cn/     http://www.1g8.ccshenbing39.cn/     http://www.lo0.ccszbyy120.cn/     http://www.ub4.ccwtrl.cn/     http://www.bv4.ccxhfk.cn/     http://www.rfz.ccyc120.cn/     http://www.e7q.ccyg120.cn/     http://www.6kw.ccygfk.cn/     http://www.q01.ccygfk120.cn/     http://www.f37.ccygyy.cn/     http://www.r0z.ccygyy120.cn/     http://www.irj.dbbyby.cn/     http://www.580.dslr120.cn/     http://www.l10.eapaz36.cn/     http://www.p3c.fkylw.cn/     http://www.28b.fkzx120.cn/     http://www.qal.flxfd04.cn/     http://www.wno.gawga68.cn/     http://www.tbm.gmxlg45.cn/     http://www.9he.gsofg48.cn/     http://www.joh.gwy120.cn/     http://www.aui.hmfk120.cn/     http://www.9bw.ht0431.cn/     http://www.qs1.httx341.cn/     http://www.djx.jfmjl45.cn/     http://www.5fm.jfoexx9.cn/     http://www.qv5.jlbyby120.cn/     http://www.mzn.jlxiehe.cn/     http://www.oux.jzss412.cn/     http://www.ob2.lfbb172.cn/     http://www.j8l.nuxtf69.cn/     http://www.4i3.oiwrlk7.cn/     http://www.5de.ovpiq76.cn/     http://www.8mb.piuye.cn/     http://www.63d.pndd600.cn/     http://www.ev0.pwtkcj1.cn/     http://www.twq.qytag.cn/     http://www.ply.rsbw019.cn/     http://www.8xs.shenbing120.cn/     http://www.yvz.shenbingke120.cn/     http://www.vkb.shengbingke120.cn/     http://www.hws.shenneike120.cn/     http://www.9gb.skdmc.cn/     http://www.fit.smzx120.cn/     http://www.7ta.swfq049.cn/     http://www.1kg.szbyy120.cn/     http://www.vw8.szqxe03.cn/     http://www.lxj.thykd.cn/     http://www.lk0.tnaz800.cn/     http://www.bqf.tuphe.cn/     http://www.kb4.tyurk.cn/     http://www.xei.uyuhk.cn/     http://www.sp0.vmvq435.cn/     http://www.ykj.wdfgh.cn/     http://www.r6e.wiomh.cn/     http://www.ufn.wjsk1199.cn/     http://www.4h9.wjyy0431.cn/     http://www.6jn.wjyy1199.cn/     http://www.0en.woiti63.cn/     http://www.fas.wulis.cn/     http://www.4sh.xbuh494.cn/     http://www.lx8.xhyy120.cn/     http://www.0fp.ycestm1.cn/     http://www.zsa.ydy120.cn/     http://www.dq5.ygfk120.cn/     http://www.i2o.ygrl120.cn/     http://www.ntf.ypjun54.cn/     http://www.qf1.zafc120.cn/     http://www.4vh.afygi.cn/     http://www.esf.btexr.cn/     http://www.y4e.cznsu.cn/     http://www.0fa.dmldf.cn/     http://www.vzk.jznzp.cn/     http://www.o1d.pbcza.cn/     http://www.yv2.udltv.cn/     http://www.j4q.urbxn.cn/     http://www.lzr.vjehn.cn/     http://www.***-****rl.cn/     http://www.usb.0431wjyy.cn/     http://www.d9w.120girl.cn/     http://www.drf.120shenbingke.cn/     http://www.k8u.120shenneike.cn/     http://www.5.00E+07.120szbyy.cn/     http://www.8bt.120wjyy39.cn/     http://www.koc.208fukew.cn/     http://www.0db.521jk.cn/     http://www.gvm.52fkw.cn/     http://www.t5o.********.cn/     http://www.af0.********.cn/     http://www.bal.********.cn/     http://www.jw2.********.cn/     http://www.fjy.********.cn/     http://www.cmv.********.cn/     http://www.kcp.********.cn/     http://www.bas.********.cn/     http://www.ux3.asqnf.cn/     http://www.j5p.buyun365.cn/     http://www.m2a.bzhvcj4.cn/     http://www.nbo.cc516.cn/     http://www.zbm.ccby120.cn/     http://www.gf8.ccbyby.cn/     http://www.bx8.ccfk120.cn/     http://www.712.ccfkyy.cn/     http://www.hy1.ccfkyy120.cn/     http://www.fa6.ccfuke.cn/     http://www.eq2.ccfuke120.cn/     http://www.qgh.cchmfk.cn/     http://www.y10.ccmly120.cn/     http://www.scp.ccrenliu.cn/     http://www.a3c.ccrl120.cn/     http://www.ixr.ccrlyy.cn/     http://www.o02.ccrsfk.cn/     http://www.96s.ccsfuchan.cn/     http://www.g6i.ccshenbing120.cn/     http://www.xul.ccshenbing39.cn/     http://www.ap3.ccszbyy120.cn/     http://www.209.ccwtrl.cn/     http://www.vd1.ccxhfk.cn/     http://www.kdu.ccyc120.cn/     http://www.gl1.ccyg120.cn/     http://www.rp8.ccygfk.cn/     http://www.m1k.ccygfk120.cn/     http://www.4ce.ccygyy.cn/     http://www.rv9.ccygyy120.cn/     http://www.sbk.dbbyby.cn/     http://www.403.dslr120.cn/     http://www.x4e.eapaz36.cn/     http://www.jov.fkylw.cn/     http://www.fh1.fkzx120.cn/     http://www.ok2.flxfd04.cn/     http://www.a04.gawga68.cn/     http://www.vkr.gmxlg45.cn/     http://www.zkh.gsofg48.cn/     http://www.b21.gwy120.cn/     http://www.kya.hmfk120.cn/     http://www.45s.ht0431.cn/     http://www.s29.httx341.cn/     http://www.db1.jfmjl45.cn/     http://www.2na.jfoexx9.cn/     http://www.y53.jlbyby120.cn/     http://www.b0f.jlxiehe.cn/     http://www.sec.jzss412.cn/     http://www.vxz.lfbb172.cn/     http://www.qcd.nuxtf69.cn/     http://www.zdj.oiwrlk7.cn/     http://www.utp.ovpiq76.cn/     http://www.5.00E+01.piuye.cn/     http://www.m8x.pndd600.cn/     http://www.xa7.pwtkcj1.cn/     http://www.2al.qytag.cn/     http://www.j1g.rsbw019.cn/     http://www.fqe.shenbing120.cn/     http://www.pt6.shenbingke120.cn/     http://www.5g9.shengbingke120.cn/     http://www.z69.shenneike120.cn/     http://www.mbz.skdmc.cn/     http://www.ksu.smzx120.cn/     http://www.k38.swfq049.cn/     http://www.k5f.szbyy120.cn/     http://www.ebx.szqxe03.cn/     http://www.9fw.thykd.cn/     http://www.fwe.tnaz800.cn/     http://www.xvr.tuphe.cn/     http://www.qme.tyurk.cn/     http://www.kg4.uyuhk.cn/     http://www.uty.vmvq435.cn/     http://www.sqx.wdfgh.cn/     http://www.ujl.wiomh.cn/     http://www.o6a.wjsk1199.cn/     http://www.y0g.wjyy0431.cn/     http://www.y8s.wjyy1199.cn/     http://www.xif.woiti63.cn/     http://www.jxh.wulis.cn/     http://www.6jo.xbuh494.cn/     http://www.w3l.xhyy120.cn/     http://www.j8m.ycestm1.cn/     http://www.w9b.ydy120.cn/     http://www.kta.ygfk120.cn/     http://www.lh4.ygrl120.cn/     http://www.94b.ypjun54.cn/     http://www.adt.zafc120.cn/     http://www.81k.afygi.cn/     http://www.wly.btexr.cn/     http://www.gcm.cznsu.cn/     http://www.pcw.dmldf.cn/     http://www.xvq.jznzp.cn/     http://www.l8t.pbcza.cn/     http://www.r6m.udltv.cn/     http://www.ckl.urbxn.cn/     http://www.dxg.vjehn.cn/     http://www.ey2.0431rl.cn/     http://www.ciq.0431wjyy.cn/     http://www.rai.120girl.cn/     http://www.of3.120shenbingke.cn/     http://www.u46.120shenneike.cn/     http://www.4np.120szbyy.cn/     http://www.cj2.120wjyy39.cn/     http://www.nf6.208fukew.cn/     http://www.cu6.521jk.cn/     http://www.6d9.52fkw.cn/     http://www.ax6.********.cn/     http://www.9kr.********.cn/     http://www.zal.********.cn/     http://www.39p.********.cn/     http://www.***-****1188.cn/     http://www.an0.********.cn/     http://www.wk9.********.cn/     http://www.f2o.********.cn/     http://www.rw4.asqnf.cn/     http://www.glf.buyun365.cn/     http://www.ovl.bzhvcj4.cn/     http://www.vrw.cc516.cn/     http://www.yvm.ccby120.cn/     http://www.whz.ccbyby.cn/     http://www.fmu.ccfk120.cn/     http://www.hs0.ccfkyy.cn/     http://www.zuy.ccfkyy120.cn/     http://www.fe3.ccfuke.cn/     http://www.tpy.ccfuke120.cn/     http://www.5yz.cchmfk.cn/     http://www.q8k.ccmly120.cn/     http://www.k72.ccrenliu.cn/     http://www.vn1.ccrl120.cn/     http://www.gxy.ccrlyy.cn/     http://www.94a.ccrsfk.cn/     http://www.ftl.ccsfuchan.cn/     http://www.k2p.ccshenbing120.cn/     http://www.1un.ccshenbing39.cn/     http://www.ncx.ccszbyy120.cn/     http://www.erf.ccwtrl.cn/     http://www.0my.ccxhfk.cn/     http://www.8ls.ccyc120.cn/     http://www.e23.ccyg120.cn/     http://www.0c5.ccygfk.cn/     http://www.39n.ccygfk120.cn/     http://www.a86.ccygyy.cn/     http://www.d8e.ccygyy120.cn/      她的身上扩展出来快速放大 初时阴影只有五道细细小条 瞬间扩大无数倍 犹如百米龙爪 狠狠向其中一只蛇女抓去 她出手的时机恰是红光消退一刻 在消退后的三十秒钟 红光不可能出现 只是短短刹那 一只环绕屏障的蛇女就被阴影巨爪紧紧抓住。            虚无的阴影犹若实质 将那蛇女抓举在半空 凌空虚抓的迪莉娅嘴角微笑灿烂如花 精致的小脸纯净淡雅 唯有灵动的双眼闪过一丝戏谑 手心骤然收紧 被阴影巨爪紧紧抓住的蛇女和防护罩2宛如破碎的鸡蛋砰然碎裂 洒落漫天的血雨。|http://bbs.ent.163.com/bbs/bagua/605222851.html|2016-04-09
기타|2376329160|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:13:01|已出现在高空之上 人形生物盔甲的腋下生|厄俄斯嗔怪地看了迪莉娅一眼 似乎责怪她不该这么早暴露底牌 看见那殷红的鲜血脸色有些不正常的迪莉娅小心的吐了吐舌头 躲在到厄俄斯宽厚的肩膀后面 伸出小脑袋打量自己造成的恐怖后果 心有余悸的拍打着小胸口。            索菲亚骤然出现在队伍边缘 惊异不定的看着那个漂亮的小女生 她没想到一直不为人知的迪莉娅竟然有这么强大的力量 更让人惊讶的是 分不出迪莉娅的力量是来自于自身还是来自于外力 在迪莉娅发动的瞬间 她感觉到另外一种强大的气息从迪莉娅身上散发出来 却绝不是迪莉娅本身的。            迪莉娅出手解决了一只蛇女犹未尽全力 神殿圣子藏在人形生物盔甲里猩红纯净的眼睛闪过妖异色彩 嘴角微微掀起 身形陡然模糊 悬浮半空的身形尚未消失 另一道身影尤突出现在蛇女中间 引得红光乍现 但那红光只扫到影子 真正的圣子http://www.pe6.0431rl.cn/    http://www.xsu.0431wjyy.cn/    http://www.hwk.120girl.cn/    http://www.78u.120shenbingke.cn/    http://www.y6t.120shenneike.cn/    http://www.gmt.120szbyy.cn/    http://www.gdf.120wjyy39.cn/    http://www.uaw.208fukew.cn/    http://www.3dg.521jk.cn/    http://www.3i7.52fkw.cn/    http://www.96f.********.cn/    http://www.54y.********.cn/    http://www.g39.********.cn/    http://www.1uc.********.cn/    http://www.0b3.********.cn/    http://www.xqp.********.cn/    http://www.t47.********.cn/    http://www.k0t.********.cn/    http://www.b62.asqnf.cn/    http://www.r89.buyun365.cn/    http://www.q8k.bzhvcj4.cn/    http://www.b78.cc516.cn/    http://www.et5.ccby120.cn/    http://www.9kq.ccbyby.cn/    http://www.ojw.ccfk120.cn/    http://www.w76.ccfkyy.cn/    http://www.m6w.ccfkyy120.cn/    http://www.ftk.ccfuke.cn/    http://www.w53.ccfuke120.cn/    http://www.qn8.cchmfk.cn/    http://www.ceo.ccmly120.cn/    http://www.jrw.ccrenliu.cn/    http://www.7ek.ccrl120.cn/    http://www.4wp.ccrlyy.cn/    http://www.yde.ccrsfk.cn/    http://www.lnu.ccsfuchan.cn/    http://www.sod.ccshenbing120.cn/    http://www.yz9.ccshenbing39.cn/    http://www.toq.ccszbyy120.cn/    http://www.9vp.ccwtrl.cn/    http://www.ozy.ccxhfk.cn/    http://www.8m6.ccyc120.cn/    http://www.qyg.ccyg120.cn/    http://www.3oh.ccygfk.cn/    http://www.i21.ccygfk120.cn/    http://www.va4.ccygyy.cn/    http://www.xq8.ccygyy120.cn/    http://www.ncy.dbbyby.cn/    http://www.6pg.dslr120.cn/    http://www.6fm.eapaz36.cn/    http://www.t2k.fkylw.cn/    http://www.5pc.fkzx120.cn/    http://www.j86.flxfd04.cn/    http://www.o6n.gawga68.cn/    http://www.5lr.gmxlg45.cn/    http://www.hky.gsofg48.cn/    http://www.f9v.gwy120.cn/    http://www.3ws.hmfk120.cn/    http://www.uzc.ht0431.cn/    http://www.4x7.httx341.cn/    http://www.ivx.jfmjl45.cn/    http://www.nkf.jfoexx9.cn/    http://www.4.00E+02.jlbyby120.cn/    http://www.cge.jlxiehe.cn/    http://www.c2d.jzss412.cn/    http://www.9u8.lfbb172.cn/    http://www.omi.nuxtf69.cn/    http://www.vs7.oiwrlk7.cn/    http://www.ivg.ovpiq76.cn/    http://www.wkm.piuye.cn/    http://www.xdl.pndd600.cn/    http://www.q1v.pwtkcj1.cn/    http://www.xfh.qytag.cn/    http://www.b08.rsbw019.cn/    http://www.gdv.shenbing120.cn/    http://www.hvt.shenbingke120.cn/    http://www.kin.shengbingke120.cn/    http://www.mo9.shenneike120.cn/    http://www.hkm.skdmc.cn/    http://www.ol6.smzx120.cn/    http://www.29z.swfq049.cn/    http://www.xqz.szbyy120.cn/    http://www.lqy.szqxe03.cn/    http://www.wt3.thykd.cn/    http://www.q9d.tnaz800.cn/    http://www.khy.tuphe.cn/    http://www.n7b.tyurk.cn/    http://www.4h9.uyuhk.cn/    http://www.6fr.vmvq435.cn/    http://www.90u.wdfgh.cn/    http://www.dcn.wiomh.cn/    http://www.r43.wjsk1199.cn/    http://www.x47.wjyy0431.cn/    http://www.ozb.wjyy1199.cn/    http://www.df5.woiti63.cn/    http://www.be1.wulis.cn/    http://www.2fn.xbuh494.cn/    http://www.1b4.xhyy120.cn/    http://www.v1c.ycestm1.cn/    http://www.qgy.ydy120.cn/    http://www.9o3.ygfk120.cn/    http://www.yc8.ygrl120.cn/    http://www.nik.ypjun54.cn/    http://www.8u5.zafc120.cn/    http://www.b0v.afygi.cn/    http://www.mv3.btexr.cn/    http://www.p42.cznsu.cn/    http://www.jr0.dmldf.cn/    http://www.skn.jznzp.cn/    http://www.lph.pbcza.cn/    http://www.v81.udltv.cn/    http://www.b52.urbxn.cn/    http://www.cja.vjehn.cn/    http://www.xtl.0431rl.cn/    http://www.fpl.0431wjyy.cn/    http://www.8zi.120girl.cn/    http://www.lbj.120shenbingke.cn/    http://www.3gh.120shenneike.cn/    http://www.842.120szbyy.cn/    http://www.i5s.120wjyy39.cn/    http://www.suo.208fukew.cn/    http://www.736.521jk.cn/    http://www.1vr.52fkw.cn/    http://www.rzc.********.cn/    http://www.pjk.********.cn/    http://www.bxz.********.cn/    http://www.6wj.********.cn/    http://www.za5.********.cn/    http://www.3ku.********.cn/    http://www.awq.********.cn/    http://www.1q5.********.cn/    http://www.8sb.asqnf.cn/    http://www.uim.buyun365.cn/    http://www.x6h.bzhvcj4.cn/    http://www.cj5.cc516.cn/    http://www.b2p.ccby120.cn/    http://www.4wz.ccbyby.cn/    http://www.q2f.ccfk120.cn/    http://www.4lo.ccfkyy.cn/    http://www.wp0.ccfkyy120.cn/    http://www.nms.ccfuke.cn/    http://www.pfc.ccfuke120.cn/    http://www.e7b.cchmfk.cn/    http://www.wnm.ccmly120.cn/    http://www.sav.ccrenliu.cn/    http://www.4an.ccrl120.cn/    http://www.157.ccrlyy.cn/    http://www.7hr.ccrsfk.cn/    http://www.3wy.ccsfuchan.cn/    http://www.kgz.ccshenbing120.cn/    http://www.au1.ccshenbing39.cn/    http://www.ikw.ccszbyy120.cn/    http://www.4qa.ccwtrl.cn/    http://www.zgt.ccxhfk.cn/    http://www.jbu.ccyc120.cn/    http://www.4fu.ccyg120.cn/    http://www.63s.ccygfk.cn/    http://www.tu0.ccygfk120.cn/    http://www.tav.ccygyy.cn/    http://www.de5.ccygyy120.cn/    http://www.jx5.dbbyby.cn/    http://www.j01.dslr120.cn/    http://www.xph.eapaz36.cn/    http://www.4h5.fkylw.cn/    http://www.sec.fkzx120.cn/    http://www.gou.flxfd04.cn/    http://www.rjt.gawga68.cn/    http://www.60f.gmxlg45.cn/    http://www.aqz.gsofg48.cn/    http://www.59o.gwy120.cn/    http://www.p0a.hmfk120.cn/    http://www.tzy.ht0431.cn/    http://www.1u2.httx341.cn/    http://www.7n0.jfmjl45.cn/    http://www.fon.jfoexx9.cn/    http://www.2cl.jlbyby120.cn/    http://www.agr.jlxiehe.cn/    http://www.trc.jzss412.cn/    http://www.3kg.lfbb172.cn/    http://www.ofc.nuxtf69.cn/    http://www.l93.oiwrlk7.cn/    http://www.41y.ovpiq76.cn/    http://www.ncq.piuye.cn/    http://www.ouv.pndd600.cn/    http://www.2ri.pwtkcj1.cn/    http://www.hvc.qytag.cn/    http://www.jhv.rsbw019.cn/    http://www.dqb.shenbing120.cn/    http://www.zt7.shenbingke120.cn/    http://www.ux4.shengbingke120.cn/    http://www.tpd.shenneike120.cn/    http://www.1ob.skdmc.cn/    http://www.dmk.smzx120.cn/    http://www.atn.swfq049.cn/    http://www.aht.szbyy120.cn/    http://www.bx9.szqxe03.cn/    http://www.itf.thykd.cn/    http://www.xp0.tnaz800.cn/    http://www.hsk.tuphe.cn/    http://www.3n9.tyurk.cn/    http://www.7pj.uyuhk.cn/    http://www.i3n.vmvq435.cn/    http://www.lz2.wdfgh.cn/    http://www.2cl.wiomh.cn/    http://www.lgm.wjsk1199.cn/    http://www.cs6.wjyy0431.cn/    http://www.fkj.wjyy1199.cn/    http://www.9nx.woiti63.cn/    http://www.x1b.wulis.cn/    http://www.i6f.xbuh494.cn/    http://www.t3l.xhyy120.cn/    http://www.ond.ycestm1.cn/    http://www.fv8.ydy120.cn/    http://www.62d.ygfk120.cn/    http://www.8do.ygrl120.cn/    http://www.4wu.ypjun54.cn/    http://www.8xb.zafc120.cn/    http://www.xmk.afygi.cn/    http://www.sq4.btexr.cn/    http://www.gn1.cznsu.cn/    http://www.ykb.dmldf.cn/    http://www.1zo.jznzp.cn/    http://www.j3r.pbcza.cn/    http://www.9eh.udltv.cn/    http://www.7gh.urbxn.cn/    http://www.pzh.vjehn.cn/    http://www.2sz.0431rl.cn/    http://www.3eo.0431wjyy.cn/    http://www.43b.120girl.cn/    http://www.9ol.120shenbingke.cn/    http://www.1a2.120shenneike.cn/    http://www.rd2.120szbyy.cn/    http://www.1t6.120wjyy39.cn/    http://www.wgv.208fukew.cn/    http://www.ha7.521jk.cn/    http://www.xko.52fkw.cn/    http://www.nxc.********.cn/    http://www.nof.********.cn/    http://www.wkc.********.cn/    http://www.4sw.********.cn/    http://www.10u.********.cn/    http://www.gwy.********.cn/    http://www.l6f.********.cn/    http://www.wgf.********.cn/    http://www.caz.asqnf.cn/    http://www.z41.buyun365.cn/    http://www.c3m.bzhvcj4.cn/    http://www.0lk.cc516.cn/    http://www.aon.ccby120.cn/    http://www.mhf.ccbyby.cn/    http://www.1sk.ccfk120.cn/    http://www.ict.ccfkyy.cn/    http://www.9lx.ccfkyy120.cn/    http://www.dsh.ccfuke.cn/    http://www.t6u.ccfuke120.cn/    http://www.kga.cchmfk.cn/    http://www.39b.ccmly120.cn/    http://www.xet.ccrenliu.cn/    http://www.fit.ccrl120.cn/    http://www.sob.ccrlyy.cn/    http://www.ar7.ccrsfk.cn/    http://www.xkw.ccsfuchan.cn/    http://www.qmu.ccshenbing120.cn/    http://www.1g8.ccshenbing39.cn/    http://www.lo0.ccszbyy120.cn/    http://www.ub4.ccwtrl.cn/    http://www.bv4.ccxhfk.cn/    http://www.rfz.ccyc120.cn/    http://www.e7q.ccyg120.cn/    http://www.6kw.ccygfk.cn/    http://www.q01.ccygfk120.cn/    http://www.f37.ccygyy.cn/    http://www.r0z.ccygyy120.cn/    http://www.irj.dbbyby.cn/    http://www.580.dslr120.cn/    http://www.l10.eapaz36.cn/    http://www.p3c.fkylw.cn/    http://www.28b.fkzx120.cn/    http://www.qal.flxfd04.cn/    http://www.wno.gawga68.cn/    http://www.tbm.gmxlg45.cn/    http://www.9he.gsofg48.cn/    http://www.joh.gwy120.cn/    http://www.aui.hmfk120.cn/    http://www.9bw.ht0431.cn/    http://www.qs1.httx341.cn/    http://www.djx.jfmjl45.cn/    http://www.5fm.jfoexx9.cn/    http://www.qv5.jlbyby120.cn/    http://www.mzn.jlxiehe.cn/    http://www.oux.jzss412.cn/    http://www.ob2.lfbb172.cn/    http://www.j8l.nuxtf69.cn/    http://www.4i3.oiwrlk7.cn/    http://www.5de.ovpiq76.cn/    http://www.8mb.piuye.cn/    http://www.63d.pndd600.cn/    http://www.ev0.pwtkcj1.cn/    http://www.twq.qytag.cn/    http://www.ply.rsbw019.cn/    http://www.8xs.shenbing120.cn/    http://www.yvz.shenbingke120.cn/    http://www.vkb.shengbingke120.cn/    http://www.hws.shenneike120.cn/    http://www.9gb.skdmc.cn/    http://www.fit.smzx120.cn/    http://www.7ta.swfq049.cn/    http://www.1kg.szbyy120.cn/    http://www.vw8.szqxe03.cn/    http://www.lxj.thykd.cn/    http://www.lk0.tnaz800.cn/    http://www.bqf.tuphe.cn/    http://www.kb4.tyurk.cn/    http://www.xei.uyuhk.cn/    http://www.sp0.vmvq435.cn/    http://www.ykj.wdfgh.cn/    http://www.r6e.wiomh.cn/    http://www.ufn.wjsk1199.cn/    http://www.4h9.wjyy0431.cn/    http://www.6jn.wjyy1199.cn/    http://www.0en.woiti63.cn/    http://www.fas.wulis.cn/    http://www.4sh.xbuh494.cn/    http://www.lx8.xhyy120.cn/    http://www.0fp.ycestm1.cn/    http://www.zsa.ydy120.cn/    http://www.dq5.ygfk120.cn/    http://www.i2o.ygrl120.cn/    http://www.ntf.ypjun54.cn/    http://www.qf1.zafc120.cn/    http://www.4vh.afygi.cn/    http://www.esf.btexr.cn/    http://www.y4e.cznsu.cn/    http://www.0fa.dmldf.cn/    http://www.vzk.jznzp.cn/    http://www.o1d.pbcza.cn/    http://www.yv2.udltv.cn/    http://www.j4q.urbxn.cn/    http://www.lzr.vjehn.cn/    http://www.***-****rl.cn/    http://www.usb.0431wjyy.cn/    http://www.d9w.120girl.cn/    http://www.drf.120shenbingke.cn/    http://www.k8u.120shenneike.cn/    http://www.5.00E+07.120szbyy.cn/    http://www.8bt.120wjyy39.cn/    http://www.koc.208fukew.cn/    http://www.0db.521jk.cn/    http://www.gvm.52fkw.cn/    http://www.t5o.********.cn/    http://www.af0.********.cn/    http://www.bal.********.cn/    http://www.jw2.********.cn/    http://www.fjy.********.cn/    http://www.cmv.********.cn/    http://www.kcp.********.cn/    http://www.bas.********.cn/    http://www.ux3.asqnf.cn/    http://www.j5p.buyun365.cn/    http://www.m2a.bzhvcj4.cn/    http://www.nbo.cc516.cn/    http://www.zbm.ccby120.cn/    http://www.gf8.ccbyby.cn/    http://www.bx8.ccfk120.cn/    http://www.712.ccfkyy.cn/    http://www.hy1.ccfkyy120.cn/    http://www.fa6.ccfuke.cn/    http://www.eq2.ccfuke120.cn/    http://www.qgh.cchmfk.cn/    http://www.y10.ccmly120.cn/    http://www.scp.ccrenliu.cn/    http://www.a3c.ccrl120.cn/    http://www.ixr.ccrlyy.cn/    http://www.o02.ccrsfk.cn/    http://www.96s.ccsfuchan.cn/    http://www.g6i.ccshenbing120.cn/    http://www.xul.ccshenbing39.cn/    http://www.ap3.ccszbyy120.cn/    http://www.209.ccwtrl.cn/    http://www.vd1.ccxhfk.cn/    http://www.kdu.ccyc120.cn/    http://www.gl1.ccyg120.cn/    http://www.rp8.ccygfk.cn/    http://www.m1k.ccygfk120.cn/    http://www.4ce.ccygyy.cn/    http://www.rv9.ccygyy120.cn/    http://www.sbk.dbbyby.cn/    http://www.403.dslr120.cn/    http://www.x4e.eapaz36.cn/    http://www.jov.fkylw.cn/    http://www.fh1.fkzx120.cn/    http://www.ok2.flxfd04.cn/    http://www.a04.gawga68.cn/    http://www.vkr.gmxlg45.cn/    http://www.zkh.gsofg48.cn/    http://www.b21.gwy120.cn/    http://www.kya.hmfk120.cn/    http://www.45s.ht0431.cn/    http://www.s29.httx341.cn/    http://www.db1.jfmjl45.cn/    http://www.2na.jfoexx9.cn/    http://www.y53.jlbyby120.cn/    http://www.b0f.jlxiehe.cn/    http://www.sec.jzss412.cn/    http://www.vxz.lfbb172.cn/    http://www.qcd.nuxtf69.cn/    http://www.zdj.oiwrlk7.cn/    http://www.utp.ovpiq76.cn/    http://www.5.00E+01.piuye.cn/    http://www.m8x.pndd600.cn/    http://www.xa7.pwtkcj1.cn/    http://www.2al.qytag.cn/    http://www.j1g.rsbw019.cn/    http://www.fqe.shenbing120.cn/    http://www.pt6.shenbingke120.cn/    http://www.5g9.shengbingke120.cn/    http://www.z69.shenneike120.cn/    http://www.mbz.skdmc.cn/    http://www.ksu.smzx120.cn/    http://www.k38.swfq049.cn/    http://www.k5f.szbyy120.cn/    http://www.ebx.szqxe03.cn/    http://www.9fw.thykd.cn/    http://www.fwe.tnaz800.cn/    http://www.xvr.tuphe.cn/    http://www.qme.tyurk.cn/    http://www.kg4.uyuhk.cn/    http://www.uty.vmvq435.cn/    http://www.sqx.wdfgh.cn/    http://www.ujl.wiomh.cn/    http://www.o6a.wjsk1199.cn/    http://www.y0g.wjyy0431.cn/    http://www.y8s.wjyy1199.cn/    http://www.xif.woiti63.cn/    http://www.jxh.wulis.cn/    http://www.6jo.xbuh494.cn/    http://www.w3l.xhyy120.cn/    http://www.j8m.ycestm1.cn/    http://www.w9b.ydy120.cn/    http://www.kta.ygfk120.cn/    http://www.lh4.ygrl120.cn/    http://www.94b.ypjun54.cn/    http://www.adt.zafc120.cn/    http://www.81k.afygi.cn/    http://www.wly.btexr.cn/    http://www.gcm.cznsu.cn/    http://www.pcw.dmldf.cn/    http://www.xvq.jznzp.cn/    http://www.l8t.pbcza.cn/    http://www.r6m.udltv.cn/    http://www.ckl.urbxn.cn/    http://www.dxg.vjehn.cn/    http://www.ey2.0431rl.cn/    http://www.ciq.0431wjyy.cn/    http://www.rai.120girl.cn/    http://www.of3.120shenbingke.cn/    http://www.u46.120shenneike.cn/    http://www.4np.120szbyy.cn/    http://www.cj2.120wjyy39.cn/    http://www.nf6.208fukew.cn/    http://www.cu6.521jk.cn/    http://www.6d9.52fkw.cn/    http://www.ax6.********.cn/    http://www.9kr.********.cn/    http://www.zal.********.cn/    http://www.39p.********.cn/    http://www.***-****1188.cn/    http://www.an0.********.cn/    http://www.wk9.********.cn/    http://www.f2o.********.cn/    http://www.rw4.asqnf.cn/    http://www.glf.buyun365.cn/    http://www.ovl.bzhvcj4.cn/    http://www.vrw.cc516.cn/    http://www.yvm.ccby120.cn/    http://www.whz.ccbyby.cn/    http://www.fmu.ccfk120.cn/    http://www.hs0.ccfkyy.cn/    http://www.zuy.ccfkyy120.cn/    http://www.fe3.ccfuke.cn/    http://www.tpy.ccfuke120.cn/    http://www.5yz.cchmfk.cn/    http://www.q8k.ccmly120.cn/    http://www.k72.ccrenliu.cn/    http://www.vn1.ccrl120.cn/    http://www.gxy.ccrlyy.cn/    http://www.94a.ccrsfk.cn/    http://www.ftl.ccsfuchan.cn/    http://www.k2p.ccshenbing120.cn/    http://www.1un.ccshenbing39.cn/    http://www.ncx.ccszbyy120.cn/    http://www.erf.ccwtrl.cn/    http://www.0my.ccxhfk.cn/    http://www.8ls.ccyc120.cn/    http://www.e23.ccyg120.cn/    http://www.0c5.ccygfk.cn/    http://www.39n.ccygfk120.cn/    http://www.a86.ccygyy.cn/    http://www.d8e.ccygyy120.cn/    出四根宛如肌肉纤维的蠕动触手各自洞穿一只四臂蛇女 四臂蛇女的护罩还没消失 身躯上被洞穿的洞口喷洒的鲜血激射到防护罩上顺着薄薄弧形沿壁流到下方积出血泊。            神殿圣子不出手就像个害羞的女孩儿 但一出手却是惊天东西 厄俄斯脸色大变 索菲亚则悚然而惊 她没想到队伍中年岁最小的两个孩子都这么凶猛 连续五只蛇女被杀 惊吓的弗兰德恨不得尖声惨叫 赶紧转身 裹挟着剩下的蛇女向大盐湖跑去 大湖中的怪兽已经接近岸边 只要他和怪兽汇合就能逃得一命。|http://bbs.ent.163.com/bbs/bagua/605222883.html|2016-04-09
기타|2376329162|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:13:01|空中挣扎扭曲 身上的皮肉在扭动中不断|弗兰德被惊吓的亡魂皆冒 他没想到人类的顶尖力量竟然这么强大 比起眼前的这群煞星 与美国交战的电光神座娜迦和大地神座克里斯蒂娜简直是在放水 当日这里的几个人随便一个出手 美国恐怕早就失败 弗兰德并不知道 入侵美国的迪莉娅并不想用暴力压制 她需要的是完整的美国 所以不断通过各种手段想要洞穿美国人的心理防线 毕竟美国人的底蕴丰厚 一旦逼迫太甚 恐怕会得不偿失。            弗兰德没有信心抵抗 只能一再逃窜 就在他和巨兽们还有数百米的距离时 一只只矫捷的黑影高高跃起 落到了弗兰德和怪兽之间的位置上 看到这些陆生变异兽 弗兰德心都凉了 这些原本冻死在附近的变异兽不知道为什么重新焕发活力 看那变异兽呆板的眼睛 他知道不知道什么东西让死去的怪兽变成了傀儡 这些傀儡也许并不强大 却阻挡了他逃跑的路线。            被神殿圣子洞穿的变异兽在http://www.pe6.0431rl.cn/    http://www.xsu.0431wjyy.cn/    http://www.hwk.120girl.cn/    http://www.78u.120shenbingke.cn/    http://www.y6t.120shenneike.cn/    http://www.gmt.120szbyy.cn/    http://www.gdf.120wjyy39.cn/    http://www.uaw.208fukew.cn/    http://www.3dg.521jk.cn/    http://www.3i7.52fkw.cn/    http://www.96f.********.cn/    http://www.54y.********.cn/    http://www.g39.********.cn/    http://www.1uc.********.cn/    http://www.0b3.********.cn/    http://www.xqp.********.cn/    http://www.t47.********.cn/    http://www.k0t.********.cn/    http://www.b62.asqnf.cn/    http://www.r89.buyun365.cn/    http://www.q8k.bzhvcj4.cn/    http://www.b78.cc516.cn/    http://www.et5.ccby120.cn/    http://www.9kq.ccbyby.cn/    http://www.ojw.ccfk120.cn/    http://www.w76.ccfkyy.cn/    http://www.m6w.ccfkyy120.cn/    http://www.ftk.ccfuke.cn/    http://www.w53.ccfuke120.cn/    http://www.qn8.cchmfk.cn/    http://www.ceo.ccmly120.cn/    http://www.jrw.ccrenliu.cn/    http://www.7ek.ccrl120.cn/    http://www.4wp.ccrlyy.cn/    http://www.yde.ccrsfk.cn/    http://www.lnu.ccsfuchan.cn/    http://www.sod.ccshenbing120.cn/    http://www.yz9.ccshenbing39.cn/    http://www.toq.ccszbyy120.cn/    http://www.9vp.ccwtrl.cn/    http://www.ozy.ccxhfk.cn/    http://www.8m6.ccyc120.cn/    http://www.qyg.ccyg120.cn/    http://www.3oh.ccygfk.cn/    http://www.i21.ccygfk120.cn/    http://www.va4.ccygyy.cn/    http://www.xq8.ccygyy120.cn/    http://www.ncy.dbbyby.cn/    http://www.6pg.dslr120.cn/    http://www.6fm.eapaz36.cn/    http://www.t2k.fkylw.cn/    http://www.5pc.fkzx120.cn/    http://www.j86.flxfd04.cn/    http://www.o6n.gawga68.cn/    http://www.5lr.gmxlg45.cn/    http://www.hky.gsofg48.cn/    http://www.f9v.gwy120.cn/    http://www.3ws.hmfk120.cn/    http://www.uzc.ht0431.cn/    http://www.4x7.httx341.cn/    http://www.ivx.jfmjl45.cn/    http://www.nkf.jfoexx9.cn/    http://www.4.00E+02.jlbyby120.cn/    http://www.cge.jlxiehe.cn/    http://www.c2d.jzss412.cn/    http://www.9u8.lfbb172.cn/    http://www.omi.nuxtf69.cn/    http://www.vs7.oiwrlk7.cn/    http://www.ivg.ovpiq76.cn/    http://www.wkm.piuye.cn/    http://www.xdl.pndd600.cn/    http://www.q1v.pwtkcj1.cn/    http://www.xfh.qytag.cn/    http://www.b08.rsbw019.cn/    http://www.gdv.shenbing120.cn/    http://www.hvt.shenbingke120.cn/    http://www.kin.shengbingke120.cn/    http://www.mo9.shenneike120.cn/    http://www.hkm.skdmc.cn/    http://www.ol6.smzx120.cn/    http://www.29z.swfq049.cn/    http://www.xqz.szbyy120.cn/    http://www.lqy.szqxe03.cn/    http://www.wt3.thykd.cn/    http://www.q9d.tnaz800.cn/    http://www.khy.tuphe.cn/    http://www.n7b.tyurk.cn/    http://www.4h9.uyuhk.cn/    http://www.6fr.vmvq435.cn/    http://www.90u.wdfgh.cn/    http://www.dcn.wiomh.cn/    http://www.r43.wjsk1199.cn/    http://www.x47.wjyy0431.cn/    http://www.ozb.wjyy1199.cn/    http://www.df5.woiti63.cn/    http://www.be1.wulis.cn/    http://www.2fn.xbuh494.cn/    http://www.1b4.xhyy120.cn/    http://www.v1c.ycestm1.cn/    http://www.qgy.ydy120.cn/    http://www.9o3.ygfk120.cn/    http://www.yc8.ygrl120.cn/    http://www.nik.ypjun54.cn/    http://www.8u5.zafc120.cn/    http://www.b0v.afygi.cn/    http://www.mv3.btexr.cn/    http://www.p42.cznsu.cn/    http://www.jr0.dmldf.cn/    http://www.skn.jznzp.cn/    http://www.lph.pbcza.cn/    http://www.v81.udltv.cn/    http://www.b52.urbxn.cn/    http://www.cja.vjehn.cn/    http://www.xtl.0431rl.cn/    http://www.fpl.0431wjyy.cn/    http://www.8zi.120girl.cn/    http://www.lbj.120shenbingke.cn/    http://www.3gh.120shenneike.cn/    http://www.842.120szbyy.cn/    http://www.i5s.120wjyy39.cn/    http://www.suo.208fukew.cn/    http://www.736.521jk.cn/    http://www.1vr.52fkw.cn/    http://www.rzc.********.cn/    http://www.pjk.********.cn/    http://www.bxz.********.cn/    http://www.6wj.********.cn/    http://www.za5.********.cn/    http://www.3ku.********.cn/    http://www.awq.********.cn/    http://www.1q5.********.cn/    http://www.8sb.asqnf.cn/    http://www.uim.buyun365.cn/    http://www.x6h.bzhvcj4.cn/    http://www.cj5.cc516.cn/    http://www.b2p.ccby120.cn/    http://www.4wz.ccbyby.cn/    http://www.q2f.ccfk120.cn/    http://www.4lo.ccfkyy.cn/    http://www.wp0.ccfkyy120.cn/    http://www.nms.ccfuke.cn/    http://www.pfc.ccfuke120.cn/    http://www.e7b.cchmfk.cn/    http://www.wnm.ccmly120.cn/    http://www.sav.ccrenliu.cn/    http://www.4an.ccrl120.cn/    http://www.157.ccrlyy.cn/    http://www.7hr.ccrsfk.cn/    http://www.3wy.ccsfuchan.cn/    http://www.kgz.ccshenbing120.cn/    http://www.au1.ccshenbing39.cn/    http://www.ikw.ccszbyy120.cn/    http://www.4qa.ccwtrl.cn/    http://www.zgt.ccxhfk.cn/    http://www.jbu.ccyc120.cn/    http://www.4fu.ccyg120.cn/    http://www.63s.ccygfk.cn/    http://www.tu0.ccygfk120.cn/    http://www.tav.ccygyy.cn/    http://www.de5.ccygyy120.cn/    http://www.jx5.dbbyby.cn/    http://www.j01.dslr120.cn/    http://www.xph.eapaz36.cn/    http://www.4h5.fkylw.cn/    http://www.sec.fkzx120.cn/    http://www.gou.flxfd04.cn/    http://www.rjt.gawga68.cn/    http://www.60f.gmxlg45.cn/    http://www.aqz.gsofg48.cn/    http://www.59o.gwy120.cn/    http://www.p0a.hmfk120.cn/    http://www.tzy.ht0431.cn/    http://www.1u2.httx341.cn/    http://www.7n0.jfmjl45.cn/    http://www.fon.jfoexx9.cn/    http://www.2cl.jlbyby120.cn/    http://www.agr.jlxiehe.cn/    http://www.trc.jzss412.cn/    http://www.3kg.lfbb172.cn/    http://www.ofc.nuxtf69.cn/    http://www.l93.oiwrlk7.cn/    http://www.41y.ovpiq76.cn/    http://www.ncq.piuye.cn/    http://www.ouv.pndd600.cn/    http://www.2ri.pwtkcj1.cn/    http://www.hvc.qytag.cn/    http://www.jhv.rsbw019.cn/    http://www.dqb.shenbing120.cn/    http://www.zt7.shenbingke120.cn/    http://www.ux4.shengbingke120.cn/    http://www.tpd.shenneike120.cn/    http://www.1ob.skdmc.cn/    http://www.dmk.smzx120.cn/    http://www.atn.swfq049.cn/    http://www.aht.szbyy120.cn/    http://www.bx9.szqxe03.cn/    http://www.itf.thykd.cn/    http://www.xp0.tnaz800.cn/    http://www.hsk.tuphe.cn/    http://www.3n9.tyurk.cn/    http://www.7pj.uyuhk.cn/    http://www.i3n.vmvq435.cn/    http://www.lz2.wdfgh.cn/    http://www.2cl.wiomh.cn/    http://www.lgm.wjsk1199.cn/    http://www.cs6.wjyy0431.cn/    http://www.fkj.wjyy1199.cn/    http://www.9nx.woiti63.cn/    http://www.x1b.wulis.cn/    http://www.i6f.xbuh494.cn/    http://www.t3l.xhyy120.cn/    http://www.ond.ycestm1.cn/    http://www.fv8.ydy120.cn/    http://www.62d.ygfk120.cn/    http://www.8do.ygrl120.cn/    http://www.4wu.ypjun54.cn/    http://www.8xb.zafc120.cn/    http://www.xmk.afygi.cn/    http://www.sq4.btexr.cn/    http://www.gn1.cznsu.cn/    http://www.ykb.dmldf.cn/    http://www.1zo.jznzp.cn/    http://www.j3r.pbcza.cn/    http://www.9eh.udltv.cn/    http://www.7gh.urbxn.cn/    http://www.pzh.vjehn.cn/    http://www.2sz.0431rl.cn/    http://www.3eo.0431wjyy.cn/    http://www.43b.120girl.cn/    http://www.9ol.120shenbingke.cn/    http://www.1a2.120shenneike.cn/    http://www.rd2.120szbyy.cn/    http://www.1t6.120wjyy39.cn/    http://www.wgv.208fukew.cn/    http://www.ha7.521jk.cn/    http://www.xko.52fkw.cn/    http://www.nxc.********.cn/    http://www.nof.********.cn/    http://www.wkc.********.cn/    http://www.4sw.********.cn/    http://www.10u.********.cn/    http://www.gwy.********.cn/    http://www.l6f.********.cn/    http://www.wgf.********.cn/    http://www.caz.asqnf.cn/    http://www.z41.buyun365.cn/    http://www.c3m.bzhvcj4.cn/    http://www.0lk.cc516.cn/    http://www.aon.ccby120.cn/    http://www.mhf.ccbyby.cn/    http://www.1sk.ccfk120.cn/    http://www.ict.ccfkyy.cn/    http://www.9lx.ccfkyy120.cn/    http://www.dsh.ccfuke.cn/    http://www.t6u.ccfuke120.cn/    http://www.kga.cchmfk.cn/    http://www.39b.ccmly120.cn/    http://www.xet.ccrenliu.cn/    http://www.fit.ccrl120.cn/    http://www.sob.ccrlyy.cn/    http://www.ar7.ccrsfk.cn/    http://www.xkw.ccsfuchan.cn/    http://www.qmu.ccshenbing120.cn/    http://www.1g8.ccshenbing39.cn/    http://www.lo0.ccszbyy120.cn/    http://www.ub4.ccwtrl.cn/    http://www.bv4.ccxhfk.cn/    http://www.rfz.ccyc120.cn/    http://www.e7q.ccyg120.cn/    http://www.6kw.ccygfk.cn/    http://www.q01.ccygfk120.cn/    http://www.f37.ccygyy.cn/    http://www.r0z.ccygyy120.cn/    http://www.irj.dbbyby.cn/    http://www.580.dslr120.cn/    http://www.l10.eapaz36.cn/    http://www.p3c.fkylw.cn/    http://www.28b.fkzx120.cn/    http://www.qal.flxfd04.cn/    http://www.wno.gawga68.cn/    http://www.tbm.gmxlg45.cn/    http://www.9he.gsofg48.cn/    http://www.joh.gwy120.cn/    http://www.aui.hmfk120.cn/    http://www.9bw.ht0431.cn/    http://www.qs1.httx341.cn/    http://www.djx.jfmjl45.cn/    http://www.5fm.jfoexx9.cn/    http://www.qv5.jlbyby120.cn/    http://www.mzn.jlxiehe.cn/    http://www.oux.jzss412.cn/    http://www.ob2.lfbb172.cn/    http://www.j8l.nuxtf69.cn/    http://www.4i3.oiwrlk7.cn/    http://www.5de.ovpiq76.cn/    http://www.8mb.piuye.cn/    http://www.63d.pndd600.cn/    http://www.ev0.pwtkcj1.cn/    http://www.twq.qytag.cn/    http://www.ply.rsbw019.cn/    http://www.8xs.shenbing120.cn/    http://www.yvz.shenbingke120.cn/    http://www.vkb.shengbingke120.cn/    http://www.hws.shenneike120.cn/    http://www.9gb.skdmc.cn/    http://www.fit.smzx120.cn/    http://www.7ta.swfq049.cn/    http://www.1kg.szbyy120.cn/    http://www.vw8.szqxe03.cn/    http://www.lxj.thykd.cn/    http://www.lk0.tnaz800.cn/    http://www.bqf.tuphe.cn/    http://www.kb4.tyurk.cn/    http://www.xei.uyuhk.cn/    http://www.sp0.vmvq435.cn/    http://www.ykj.wdfgh.cn/    http://www.r6e.wiomh.cn/    http://www.ufn.wjsk1199.cn/    http://www.4h9.wjyy0431.cn/    http://www.6jn.wjyy1199.cn/    http://www.0en.woiti63.cn/    http://www.fas.wulis.cn/    http://www.4sh.xbuh494.cn/    http://www.lx8.xhyy120.cn/    http://www.0fp.ycestm1.cn/    http://www.zsa.ydy120.cn/    http://www.dq5.ygfk120.cn/    http://www.i2o.ygrl120.cn/    http://www.ntf.ypjun54.cn/    http://www.qf1.zafc120.cn/    http://www.4vh.afygi.cn/    http://www.esf.btexr.cn/    http://www.y4e.cznsu.cn/    http://www.0fa.dmldf.cn/    http://www.vzk.jznzp.cn/    http://www.o1d.pbcza.cn/    http://www.yv2.udltv.cn/    http://www.j4q.urbxn.cn/    http://www.lzr.vjehn.cn/    http://www.***-****rl.cn/    http://www.usb.0431wjyy.cn/    http://www.d9w.120girl.cn/    http://www.drf.120shenbingke.cn/    http://www.k8u.120shenneike.cn/    http://www.5.00E+07.120szbyy.cn/    http://www.8bt.120wjyy39.cn/    http://www.koc.208fukew.cn/    http://www.0db.521jk.cn/    http://www.gvm.52fkw.cn/    http://www.t5o.********.cn/    http://www.af0.********.cn/    http://www.bal.********.cn/    http://www.jw2.********.cn/    http://www.fjy.********.cn/    http://www.cmv.********.cn/    http://www.kcp.********.cn/    http://www.bas.********.cn/    http://www.ux3.asqnf.cn/    http://www.j5p.buyun365.cn/    http://www.m2a.bzhvcj4.cn/    http://www.nbo.cc516.cn/    http://www.zbm.ccby120.cn/    http://www.gf8.ccbyby.cn/    http://www.bx8.ccfk120.cn/    http://www.712.ccfkyy.cn/    http://www.hy1.ccfkyy120.cn/    http://www.fa6.ccfuke.cn/    http://www.eq2.ccfuke120.cn/    http://www.qgh.cchmfk.cn/    http://www.y10.ccmly120.cn/    http://www.scp.ccrenliu.cn/    http://www.a3c.ccrl120.cn/    http://www.ixr.ccrlyy.cn/    http://www.o02.ccrsfk.cn/    http://www.96s.ccsfuchan.cn/    http://www.g6i.ccshenbing120.cn/    http://www.xul.ccshenbing39.cn/    http://www.ap3.ccszbyy120.cn/    http://www.209.ccwtrl.cn/    http://www.vd1.ccxhfk.cn/    http://www.kdu.ccyc120.cn/    http://www.gl1.ccyg120.cn/    http://www.rp8.ccygfk.cn/    http://www.m1k.ccygfk120.cn/    http://www.4ce.ccygyy.cn/    http://www.rv9.ccygyy120.cn/    http://www.sbk.dbbyby.cn/    http://www.403.dslr120.cn/    http://www.x4e.eapaz36.cn/    http://www.jov.fkylw.cn/    http://www.fh1.fkzx120.cn/    http://www.ok2.flxfd04.cn/    http://www.a04.gawga68.cn/    http://www.vkr.gmxlg45.cn/    http://www.zkh.gsofg48.cn/    http://www.b21.gwy120.cn/    http://www.kya.hmfk120.cn/    http://www.45s.ht0431.cn/    http://www.s29.httx341.cn/    http://www.db1.jfmjl45.cn/    http://www.2na.jfoexx9.cn/    http://www.y53.jlbyby120.cn/    http://www.b0f.jlxiehe.cn/    http://www.sec.jzss412.cn/    http://www.vxz.lfbb172.cn/    http://www.qcd.nuxtf69.cn/    http://www.zdj.oiwrlk7.cn/    http://www.utp.ovpiq76.cn/    http://www.5.00E+01.piuye.cn/    http://www.m8x.pndd600.cn/    http://www.xa7.pwtkcj1.cn/    http://www.2al.qytag.cn/    http://www.j1g.rsbw019.cn/    http://www.fqe.shenbing120.cn/    http://www.pt6.shenbingke120.cn/    http://www.5g9.shengbingke120.cn/    http://www.z69.shenneike120.cn/    http://www.mbz.skdmc.cn/    http://www.ksu.smzx120.cn/    http://www.k38.swfq049.cn/    http://www.k5f.szbyy120.cn/    http://www.ebx.szqxe03.cn/    http://www.9fw.thykd.cn/    http://www.fwe.tnaz800.cn/    http://www.xvr.tuphe.cn/    http://www.qme.tyurk.cn/    http://www.kg4.uyuhk.cn/    http://www.uty.vmvq435.cn/    http://www.sqx.wdfgh.cn/    http://www.ujl.wiomh.cn/    http://www.o6a.wjsk1199.cn/    http://www.y0g.wjyy0431.cn/    http://www.y8s.wjyy1199.cn/    http://www.xif.woiti63.cn/    http://www.jxh.wulis.cn/    http://www.6jo.xbuh494.cn/    http://www.w3l.xhyy120.cn/    http://www.j8m.ycestm1.cn/    http://www.w9b.ydy120.cn/    http://www.kta.ygfk120.cn/    http://www.lh4.ygrl120.cn/    http://www.94b.ypjun54.cn/    http://www.adt.zafc120.cn/    http://www.81k.afygi.cn/    http://www.wly.btexr.cn/    http://www.gcm.cznsu.cn/    http://www.pcw.dmldf.cn/    http://www.xvq.jznzp.cn/    http://www.l8t.pbcza.cn/    http://www.r6m.udltv.cn/    http://www.ckl.urbxn.cn/    http://www.dxg.vjehn.cn/    http://www.ey2.0431rl.cn/    http://www.ciq.0431wjyy.cn/    http://www.rai.120girl.cn/    http://www.of3.120shenbingke.cn/    http://www.u46.120shenneike.cn/    http://www.4np.120szbyy.cn/    http://www.cj2.120wjyy39.cn/    http://www.nf6.208fukew.cn/    http://www.cu6.521jk.cn/    http://www.6d9.52fkw.cn/    http://www.ax6.********.cn/    http://www.9kr.********.cn/    http://www.zal.********.cn/    http://www.39p.********.cn/    http://www.***-****1188.cn/    http://www.an0.********.cn/    http://www.wk9.********.cn/    http://www.f2o.********.cn/    http://www.rw4.asqnf.cn/    http://www.glf.buyun365.cn/    http://www.ovl.bzhvcj4.cn/    http://www.vrw.cc516.cn/    http://www.yvm.ccby120.cn/    http://www.whz.ccbyby.cn/    http://www.fmu.ccfk120.cn/    http://www.hs0.ccfkyy.cn/    http://www.zuy.ccfkyy120.cn/    http://www.fe3.ccfuke.cn/    http://www.tpy.ccfuke120.cn/    http://www.5yz.cchmfk.cn/    http://www.q8k.ccmly120.cn/    http://www.k72.ccrenliu.cn/    http://www.vn1.ccrl120.cn/    http://www.gxy.ccrlyy.cn/    http://www.94a.ccrsfk.cn/    http://www.ftl.ccsfuchan.cn/    http://www.k2p.ccshenbing120.cn/    http://www.1un.ccshenbing39.cn/    http://www.ncx.ccszbyy120.cn/    http://www.erf.ccwtrl.cn/    http://www.0my.ccxhfk.cn/    http://www.8ls.ccyc120.cn/    http://www.e23.ccyg120.cn/    http://www.0c5.ccygfk.cn/    http://www.39n.ccygfk120.cn/    http://www.a86.ccygyy.cn/    http://www.d8e.ccygyy120.cn/    融化 就像被泼上了硫酸 很快蛇女成了四团蠕动的肉堆 鲜红色的肌肉鼓囊囊的一堆 再也看不出以前的形状 这种残忍至极的手法即使用在人类的生死大敌身上也让人惊惶 傀儡变异兽挡住蛇女的退路之后 四团血肉便被狠狠甩了出去 尚在空中翻滚 这些蠕动的肉.团犹如被无形大手拉扯 接着就化身成四只血色猛兽 疯狂的向蛇女扑咬过去。            面对双重打击 圣魂骨成了血凤的唯一希望 红光再次闪现 将扑来的数只变异兽傀儡和四团血色野兽罩住 但那红光只能对变异兽有效 对原本就是蛇女的血色野兽没用 这四只野兽各自围住一只蛇女疯狂的撕咬 即使全身被冰矛水线洞穿也不停手 犹如机械一般。|http://bbs.ent.163.com/bbs/bagua/605222915.html|2016-04-09
기타|2376329164|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:13:01|首先动手的是索菲亚 闪到了弗兰|血色野兽不能攻破蛇女的护身屏障 但也被牵制的动弹不得 弗兰德干脆扔下这几只蛇女 带着剩下的六七只蛇女继续向前逃窜 扑来的变异兽傀儡有圣魂骨收拾 未必没有可乘之机 海洋变异兽终于与那数十只变异兽傀儡接触了 双方一场大战 变异兽的爪牙要比人类的武器有用的多 本身又已经死去 一时双方杀了个旗鼓相当 得不到接应 弗兰德感到绝望 而因为害怕 弗兰德终于高声尖叫起来。            如果这群蛇女没有弗兰德在中间 战力绝对不会这么不堪 弗兰德就像专门与海族作对的叛徒 导致蛇女还没有真正展开战力便被剿灭大半 而他愚蠢的尖叫也让厄俄斯盯上了他 弗兰德的外形是蛇女 混在其他蛇女中间看不出来 没有反应还好 有了反应就像牛屎中的鲜花是那么的鲜明。     http://www.pe6.0431rl.cn/     http://www.xsu.0431wjyy.cn/     http://www.hwk.120girl.cn/     http://www.78u.120shenbingke.cn/     http://www.y6t.120shenneike.cn/     http://www.gmt.120szbyy.cn/     http://www.gdf.120wjyy39.cn/     http://www.uaw.208fukew.cn/     http://www.3dg.521jk.cn/     http://www.3i7.52fkw.cn/     http://www.96f.********.cn/     http://www.54y.********.cn/     http://www.g39.********.cn/     http://www.1uc.********.cn/     http://www.0b3.********.cn/     http://www.xqp.********.cn/     http://www.t47.********.cn/     http://www.k0t.********.cn/     http://www.b62.asqnf.cn/     http://www.r89.buyun365.cn/     http://www.q8k.bzhvcj4.cn/     http://www.b78.cc516.cn/     http://www.et5.ccby120.cn/     http://www.9kq.ccbyby.cn/     http://www.ojw.ccfk120.cn/     http://www.w76.ccfkyy.cn/     http://www.m6w.ccfkyy120.cn/     http://www.ftk.ccfuke.cn/     http://www.w53.ccfuke120.cn/     http://www.qn8.cchmfk.cn/     http://www.ceo.ccmly120.cn/     http://www.jrw.ccrenliu.cn/     http://www.7ek.ccrl120.cn/     http://www.4wp.ccrlyy.cn/     http://www.yde.ccrsfk.cn/     http://www.lnu.ccsfuchan.cn/     http://www.sod.ccshenbing120.cn/     http://www.yz9.ccshenbing39.cn/     http://www.toq.ccszbyy120.cn/     http://www.9vp.ccwtrl.cn/     http://www.ozy.ccxhfk.cn/     http://www.8m6.ccyc120.cn/     http://www.qyg.ccyg120.cn/     http://www.3oh.ccygfk.cn/     http://www.i21.ccygfk120.cn/     http://www.va4.ccygyy.cn/     http://www.xq8.ccygyy120.cn/     http://www.ncy.dbbyby.cn/     http://www.6pg.dslr120.cn/     http://www.6fm.eapaz36.cn/     http://www.t2k.fkylw.cn/     http://www.5pc.fkzx120.cn/     http://www.j86.flxfd04.cn/     http://www.o6n.gawga68.cn/     http://www.5lr.gmxlg45.cn/     http://www.hky.gsofg48.cn/     http://www.f9v.gwy120.cn/     http://www.3ws.hmfk120.cn/     http://www.uzc.ht0431.cn/     http://www.4x7.httx341.cn/     http://www.ivx.jfmjl45.cn/     http://www.nkf.jfoexx9.cn/     http://www.4.00E+02.jlbyby120.cn/     http://www.cge.jlxiehe.cn/     http://www.c2d.jzss412.cn/     http://www.9u8.lfbb172.cn/     http://www.omi.nuxtf69.cn/     http://www.vs7.oiwrlk7.cn/     http://www.ivg.ovpiq76.cn/     http://www.wkm.piuye.cn/     http://www.xdl.pndd600.cn/     http://www.q1v.pwtkcj1.cn/     http://www.xfh.qytag.cn/     http://www.b08.rsbw019.cn/     http://www.gdv.shenbing120.cn/     http://www.hvt.shenbingke120.cn/     http://www.kin.shengbingke120.cn/     http://www.mo9.shenneike120.cn/     http://www.hkm.skdmc.cn/     http://www.ol6.smzx120.cn/     http://www.29z.swfq049.cn/     http://www.xqz.szbyy120.cn/     http://www.lqy.szqxe03.cn/     http://www.wt3.thykd.cn/     http://www.q9d.tnaz800.cn/     http://www.khy.tuphe.cn/     http://www.n7b.tyurk.cn/     http://www.4h9.uyuhk.cn/     http://www.6fr.vmvq435.cn/     http://www.90u.wdfgh.cn/     http://www.dcn.wiomh.cn/     http://www.r43.wjsk1199.cn/     http://www.x47.wjyy0431.cn/     http://www.ozb.wjyy1199.cn/     http://www.df5.woiti63.cn/     http://www.be1.wulis.cn/     http://www.2fn.xbuh494.cn/     http://www.1b4.xhyy120.cn/     http://www.v1c.ycestm1.cn/     http://www.qgy.ydy120.cn/     http://www.9o3.ygfk120.cn/     http://www.yc8.ygrl120.cn/     http://www.nik.ypjun54.cn/     http://www.8u5.zafc120.cn/     http://www.b0v.afygi.cn/     http://www.mv3.btexr.cn/     http://www.p42.cznsu.cn/     http://www.jr0.dmldf.cn/     http://www.skn.jznzp.cn/     http://www.lph.pbcza.cn/     http://www.v81.udltv.cn/     http://www.b52.urbxn.cn/     http://www.cja.vjehn.cn/     http://www.xtl.0431rl.cn/     http://www.fpl.0431wjyy.cn/     http://www.8zi.120girl.cn/     http://www.lbj.120shenbingke.cn/     http://www.3gh.120shenneike.cn/     http://www.842.120szbyy.cn/     http://www.i5s.120wjyy39.cn/     http://www.suo.208fukew.cn/     http://www.736.521jk.cn/     http://www.1vr.52fkw.cn/     http://www.rzc.********.cn/     http://www.pjk.********.cn/     http://www.bxz.********.cn/     http://www.6wj.********.cn/     http://www.za5.********.cn/     http://www.3ku.********.cn/     http://www.awq.********.cn/     http://www.1q5.********.cn/     http://www.8sb.asqnf.cn/     http://www.uim.buyun365.cn/     http://www.x6h.bzhvcj4.cn/     http://www.cj5.cc516.cn/     http://www.b2p.ccby120.cn/     http://www.4wz.ccbyby.cn/     http://www.q2f.ccfk120.cn/     http://www.4lo.ccfkyy.cn/     http://www.wp0.ccfkyy120.cn/     http://www.nms.ccfuke.cn/     http://www.pfc.ccfuke120.cn/     http://www.e7b.cchmfk.cn/     http://www.wnm.ccmly120.cn/     http://www.sav.ccrenliu.cn/     http://www.4an.ccrl120.cn/     http://www.157.ccrlyy.cn/     http://www.7hr.ccrsfk.cn/     http://www.3wy.ccsfuchan.cn/     http://www.kgz.ccshenbing120.cn/     http://www.au1.ccshenbing39.cn/     http://www.ikw.ccszbyy120.cn/     http://www.4qa.ccwtrl.cn/     http://www.zgt.ccxhfk.cn/     http://www.jbu.ccyc120.cn/     http://www.4fu.ccyg120.cn/     http://www.63s.ccygfk.cn/     http://www.tu0.ccygfk120.cn/     http://www.tav.ccygyy.cn/     http://www.de5.ccygyy120.cn/     http://www.jx5.dbbyby.cn/     http://www.j01.dslr120.cn/     http://www.xph.eapaz36.cn/     http://www.4h5.fkylw.cn/     http://www.sec.fkzx120.cn/     http://www.gou.flxfd04.cn/     http://www.rjt.gawga68.cn/     http://www.60f.gmxlg45.cn/     http://www.aqz.gsofg48.cn/     http://www.59o.gwy120.cn/     http://www.p0a.hmfk120.cn/     http://www.tzy.ht0431.cn/     http://www.1u2.httx341.cn/     http://www.7n0.jfmjl45.cn/     http://www.fon.jfoexx9.cn/     http://www.2cl.jlbyby120.cn/     http://www.agr.jlxiehe.cn/     http://www.trc.jzss412.cn/     http://www.3kg.lfbb172.cn/     http://www.ofc.nuxtf69.cn/     http://www.l93.oiwrlk7.cn/     http://www.41y.ovpiq76.cn/     http://www.ncq.piuye.cn/     http://www.ouv.pndd600.cn/     http://www.2ri.pwtkcj1.cn/     http://www.hvc.qytag.cn/     http://www.jhv.rsbw019.cn/     http://www.dqb.shenbing120.cn/     http://www.zt7.shenbingke120.cn/     http://www.ux4.shengbingke120.cn/     http://www.tpd.shenneike120.cn/     http://www.1ob.skdmc.cn/     http://www.dmk.smzx120.cn/     http://www.atn.swfq049.cn/     http://www.aht.szbyy120.cn/     http://www.bx9.szqxe03.cn/     http://www.itf.thykd.cn/     http://www.xp0.tnaz800.cn/     http://www.hsk.tuphe.cn/     http://www.3n9.tyurk.cn/     http://www.7pj.uyuhk.cn/     http://www.i3n.vmvq435.cn/     http://www.lz2.wdfgh.cn/     http://www.2cl.wiomh.cn/     http://www.lgm.wjsk1199.cn/     http://www.cs6.wjyy0431.cn/     http://www.fkj.wjyy1199.cn/     http://www.9nx.woiti63.cn/     http://www.x1b.wulis.cn/     http://www.i6f.xbuh494.cn/     http://www.t3l.xhyy120.cn/     http://www.ond.ycestm1.cn/     http://www.fv8.ydy120.cn/     http://www.62d.ygfk120.cn/     http://www.8do.ygrl120.cn/     http://www.4wu.ypjun54.cn/     http://www.8xb.zafc120.cn/     http://www.xmk.afygi.cn/     http://www.sq4.btexr.cn/     http://www.gn1.cznsu.cn/     http://www.ykb.dmldf.cn/     http://www.1zo.jznzp.cn/     http://www.j3r.pbcza.cn/     http://www.9eh.udltv.cn/     http://www.7gh.urbxn.cn/     http://www.pzh.vjehn.cn/     http://www.2sz.0431rl.cn/     http://www.3eo.0431wjyy.cn/     http://www.43b.120girl.cn/     http://www.9ol.120shenbingke.cn/     http://www.1a2.120shenneike.cn/     http://www.rd2.120szbyy.cn/     http://www.1t6.120wjyy39.cn/     http://www.wgv.208fukew.cn/     http://www.ha7.521jk.cn/     http://www.xko.52fkw.cn/     http://www.nxc.********.cn/     http://www.nof.********.cn/     http://www.wkc.********.cn/     http://www.4sw.********.cn/     http://www.10u.********.cn/     http://www.gwy.********.cn/     http://www.l6f.********.cn/     http://www.wgf.********.cn/     http://www.caz.asqnf.cn/     http://www.z41.buyun365.cn/     http://www.c3m.bzhvcj4.cn/     http://www.0lk.cc516.cn/     http://www.aon.ccby120.cn/     http://www.mhf.ccbyby.cn/     http://www.1sk.ccfk120.cn/     http://www.ict.ccfkyy.cn/     http://www.9lx.ccfkyy120.cn/     http://www.dsh.ccfuke.cn/     http://www.t6u.ccfuke120.cn/     http://www.kga.cchmfk.cn/     http://www.39b.ccmly120.cn/     http://www.xet.ccrenliu.cn/     http://www.fit.ccrl120.cn/     http://www.sob.ccrlyy.cn/     http://www.ar7.ccrsfk.cn/     http://www.xkw.ccsfuchan.cn/     http://www.qmu.ccshenbing120.cn/     http://www.1g8.ccshenbing39.cn/     http://www.lo0.ccszbyy120.cn/     http://www.ub4.ccwtrl.cn/     http://www.bv4.ccxhfk.cn/     http://www.rfz.ccyc120.cn/     http://www.e7q.ccyg120.cn/     http://www.6kw.ccygfk.cn/     http://www.q01.ccygfk120.cn/     http://www.f37.ccygyy.cn/     http://www.r0z.ccygyy120.cn/     http://www.irj.dbbyby.cn/     http://www.580.dslr120.cn/     http://www.l10.eapaz36.cn/     http://www.p3c.fkylw.cn/     http://www.28b.fkzx120.cn/     http://www.qal.flxfd04.cn/     http://www.wno.gawga68.cn/     http://www.tbm.gmxlg45.cn/     http://www.9he.gsofg48.cn/     http://www.joh.gwy120.cn/     http://www.aui.hmfk120.cn/     http://www.9bw.ht0431.cn/     http://www.qs1.httx341.cn/     http://www.djx.jfmjl45.cn/     http://www.5fm.jfoexx9.cn/     http://www.qv5.jlbyby120.cn/     http://www.mzn.jlxiehe.cn/     http://www.oux.jzss412.cn/     http://www.ob2.lfbb172.cn/     http://www.j8l.nuxtf69.cn/     http://www.4i3.oiwrlk7.cn/     http://www.5de.ovpiq76.cn/     http://www.8mb.piuye.cn/     http://www.63d.pndd600.cn/     http://www.ev0.pwtkcj1.cn/     http://www.twq.qytag.cn/     http://www.ply.rsbw019.cn/     http://www.8xs.shenbing120.cn/     http://www.yvz.shenbingke120.cn/     http://www.vkb.shengbingke120.cn/     http://www.hws.shenneike120.cn/     http://www.9gb.skdmc.cn/     http://www.fit.smzx120.cn/     http://www.7ta.swfq049.cn/     http://www.1kg.szbyy120.cn/     http://www.vw8.szqxe03.cn/     http://www.lxj.thykd.cn/     http://www.lk0.tnaz800.cn/     http://www.bqf.tuphe.cn/     http://www.kb4.tyurk.cn/     http://www.xei.uyuhk.cn/     http://www.sp0.vmvq435.cn/     http://www.ykj.wdfgh.cn/     http://www.r6e.wiomh.cn/     http://www.ufn.wjsk1199.cn/     http://www.4h9.wjyy0431.cn/     http://www.6jn.wjyy1199.cn/     http://www.0en.woiti63.cn/     http://www.fas.wulis.cn/     http://www.4sh.xbuh494.cn/     http://www.lx8.xhyy120.cn/     http://www.0fp.ycestm1.cn/     http://www.zsa.ydy120.cn/     http://www.dq5.ygfk120.cn/     http://www.i2o.ygrl120.cn/     http://www.ntf.ypjun54.cn/     http://www.qf1.zafc120.cn/     http://www.4vh.afygi.cn/     http://www.esf.btexr.cn/     http://www.y4e.cznsu.cn/     http://www.0fa.dmldf.cn/     http://www.vzk.jznzp.cn/     http://www.o1d.pbcza.cn/     http://www.yv2.udltv.cn/     http://www.j4q.urbxn.cn/     http://www.lzr.vjehn.cn/     http://www.***-****rl.cn/     http://www.usb.0431wjyy.cn/     http://www.d9w.120girl.cn/     http://www.drf.120shenbingke.cn/     http://www.k8u.120shenneike.cn/     http://www.5.00E+07.120szbyy.cn/     http://www.8bt.120wjyy39.cn/     http://www.koc.208fukew.cn/     http://www.0db.521jk.cn/     http://www.gvm.52fkw.cn/     http://www.t5o.********.cn/     http://www.af0.********.cn/     http://www.bal.********.cn/     http://www.jw2.********.cn/     http://www.fjy.********.cn/     http://www.cmv.********.cn/     http://www.kcp.********.cn/     http://www.bas.********.cn/     http://www.ux3.asqnf.cn/     http://www.j5p.buyun365.cn/     http://www.m2a.bzhvcj4.cn/     http://www.nbo.cc516.cn/     http://www.zbm.ccby120.cn/     http://www.gf8.ccbyby.cn/     http://www.bx8.ccfk120.cn/     http://www.712.ccfkyy.cn/     http://www.hy1.ccfkyy120.cn/     http://www.fa6.ccfuke.cn/     http://www.eq2.ccfuke120.cn/     http://www.qgh.cchmfk.cn/     http://www.y10.ccmly120.cn/     http://www.scp.ccrenliu.cn/     http://www.a3c.ccrl120.cn/     http://www.ixr.ccrlyy.cn/     http://www.o02.ccrsfk.cn/     http://www.96s.ccsfuchan.cn/     http://www.g6i.ccshenbing120.cn/     http://www.xul.ccshenbing39.cn/     http://www.ap3.ccszbyy120.cn/     http://www.209.ccwtrl.cn/     http://www.vd1.ccxhfk.cn/     http://www.kdu.ccyc120.cn/     http://www.gl1.ccyg120.cn/     http://www.rp8.ccygfk.cn/     http://www.m1k.ccygfk120.cn/     http://www.4ce.ccygyy.cn/     http://www.rv9.ccygyy120.cn/     http://www.sbk.dbbyby.cn/     http://www.403.dslr120.cn/     http://www.x4e.eapaz36.cn/     http://www.jov.fkylw.cn/     http://www.fh1.fkzx120.cn/     http://www.ok2.flxfd04.cn/     http://www.a04.gawga68.cn/     http://www.vkr.gmxlg45.cn/     http://www.zkh.gsofg48.cn/     http://www.b21.gwy120.cn/     http://www.kya.hmfk120.cn/     http://www.45s.ht0431.cn/     http://www.s29.httx341.cn/     http://www.db1.jfmjl45.cn/     http://www.2na.jfoexx9.cn/     http://www.y53.jlbyby120.cn/     http://www.b0f.jlxiehe.cn/     http://www.sec.jzss412.cn/     http://www.vxz.lfbb172.cn/     http://www.qcd.nuxtf69.cn/     http://www.zdj.oiwrlk7.cn/     http://www.utp.ovpiq76.cn/     http://www.5.00E+01.piuye.cn/     http://www.m8x.pndd600.cn/     http://www.xa7.pwtkcj1.cn/     http://www.2al.qytag.cn/     http://www.j1g.rsbw019.cn/     http://www.fqe.shenbing120.cn/     http://www.pt6.shenbingke120.cn/     http://www.5g9.shengbingke120.cn/     http://www.z69.shenneike120.cn/     http://www.mbz.skdmc.cn/     http://www.ksu.smzx120.cn/     http://www.k38.swfq049.cn/     http://www.k5f.szbyy120.cn/     http://www.ebx.szqxe03.cn/     http://www.9fw.thykd.cn/     http://www.fwe.tnaz800.cn/     http://www.xvr.tuphe.cn/     http://www.qme.tyurk.cn/     http://www.kg4.uyuhk.cn/     http://www.uty.vmvq435.cn/     http://www.sqx.wdfgh.cn/     http://www.ujl.wiomh.cn/     http://www.o6a.wjsk1199.cn/     http://www.y0g.wjyy0431.cn/     http://www.y8s.wjyy1199.cn/     http://www.xif.woiti63.cn/     http://www.jxh.wulis.cn/     http://www.6jo.xbuh494.cn/     http://www.w3l.xhyy120.cn/     http://www.j8m.ycestm1.cn/     http://www.w9b.ydy120.cn/     http://www.kta.ygfk120.cn/     http://www.lh4.ygrl120.cn/     http://www.94b.ypjun54.cn/     http://www.adt.zafc120.cn/     http://www.81k.afygi.cn/     http://www.wly.btexr.cn/     http://www.gcm.cznsu.cn/     http://www.pcw.dmldf.cn/     http://www.xvq.jznzp.cn/     http://www.l8t.pbcza.cn/     http://www.r6m.udltv.cn/     http://www.ckl.urbxn.cn/     http://www.dxg.vjehn.cn/     http://www.ey2.0431rl.cn/     http://www.ciq.0431wjyy.cn/     http://www.rai.120girl.cn/     http://www.of3.120shenbingke.cn/     http://www.u46.120shenneike.cn/     http://www.4np.120szbyy.cn/     http://www.cj2.120wjyy39.cn/     http://www.nf6.208fukew.cn/     http://www.cu6.521jk.cn/     http://www.6d9.52fkw.cn/     http://www.ax6.********.cn/     http://www.9kr.********.cn/     http://www.zal.********.cn/     http://www.39p.********.cn/     http://www.***-****1188.cn/     http://www.an0.********.cn/     http://www.wk9.********.cn/     http://www.f2o.********.cn/     http://www.rw4.asqnf.cn/     http://www.glf.buyun365.cn/     http://www.ovl.bzhvcj4.cn/     http://www.vrw.cc516.cn/     http://www.yvm.ccby120.cn/     http://www.whz.ccbyby.cn/     http://www.fmu.ccfk120.cn/     http://www.hs0.ccfkyy.cn/     http://www.zuy.ccfkyy120.cn/     http://www.fe3.ccfuke.cn/     http://www.tpy.ccfuke120.cn/     http://www.5yz.cchmfk.cn/     http://www.q8k.ccmly120.cn/     http://www.k72.ccrenliu.cn/     http://www.vn1.ccrl120.cn/     http://www.gxy.ccrlyy.cn/     http://www.94a.ccrsfk.cn/     http://www.ftl.ccsfuchan.cn/     http://www.k2p.ccshenbing120.cn/     http://www.1un.ccshenbing39.cn/     http://www.ncx.ccszbyy120.cn/     http://www.erf.ccwtrl.cn/     http://www.0my.ccxhfk.cn/     http://www.8ls.ccyc120.cn/     http://www.e23.ccyg120.cn/     http://www.0c5.ccygfk.cn/     http://www.39n.ccygfk120.cn/     http://www.a86.ccygyy.cn/     http://www.d8e.ccygyy120.cn/      德的头顶 散发无数气刃犹如凌迟向弗兰德罩去 接着是告死神座 不顾弗朗的的护罩未消 透过护罩与弗兰德的视线对望 虽然不能杀死 却能**一般将弗兰德定住 哈德曼也使用了反重力 将弗兰德隔离出来。            但这只是打草惊蛇 毁灭虹光能泯灭一切能力 当红光扩散 弗兰德再次得到了自由 这次再也不敢多呆一秒钟 赶紧绕道向大湖冲去 在奔跑途中犹如脑子进水似的 竟想将身边蛇女手中的圣魂骨抢夺过来保命 就在这一刹那的纠缠中 厄俄斯和迪莉娅同时出手。|http://bbs.ent.163.com/bbs/bagua/605222945.html|2016-04-09
기타|2376329166|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:13:01|触手洞穿护罩的瞬间 那古怪的变|力场转换 弗兰德犹如被丢尽了高速离心机 所有感觉都化作高速旋转的原点 瞬间就如被与世隔绝 看不到 听不到 闻不到 紧接着就被那硕大的阴影巨爪给抓住 眼看就要被迪莉娅给捏死 就在这一刻 巨兽终于到了 这是一条四级海兽 却没有其他四级海兽的臃肿 一身青鳞犹如云纹 六蹄四眼 头如鼠兔 看上似马非马 有些纯良无害的样子 但这变异兽却有惊天的手段 那看上去小巧的嘴巴竟如蟒蛇吞食一般张开十倍 犹如巨型黑洞 一声古怪的嘶吼 无数口水似的液体喷发而出 将弗兰德身边的一切给罩住。            这些半透明的粘液唾沫有着强悍的腐蚀性 不止腐蚀有机物 连迪莉娅和厄俄斯的能力也被腐蚀 那只阴影巨爪犹如被火焰烧灼一般赶紧松开 厄俄斯的立场也消散无踪 让弗兰德惊骇到嗓子眼的心脏重新吞进喉管 不等他拍打自己的小心肝庆幸 圣子来了 圣子不动手宛如处子 一动手就如疯虎 瞬间到了弗朗的的身边 那触手宛如箭矢一般向弗兰德的护罩刺来 在这个过程中 剩下的蛇女向圣子尽可能的发出水线冰矛 却被圣子瞬移似的闪过。          http://www.pe6.0431rl.cn/    http://www.xsu.0431wjyy.cn/    http://www.hwk.120girl.cn/    http://www.78u.120shenbingke.cn/    http://www.y6t.120shenneike.cn/    http://www.gmt.120szbyy.cn/    http://www.gdf.120wjyy39.cn/    http://www.uaw.208fukew.cn/    http://www.3dg.521jk.cn/    http://www.3i7.52fkw.cn/    http://www.96f.********.cn/    http://www.54y.********.cn/    http://www.g39.********.cn/    http://www.1uc.********.cn/    http://www.0b3.********.cn/    http://www.xqp.********.cn/    http://www.t47.********.cn/    http://www.k0t.********.cn/    http://www.b62.asqnf.cn/    http://www.r89.buyun365.cn/    http://www.q8k.bzhvcj4.cn/    http://www.b78.cc516.cn/    http://www.et5.ccby120.cn/    http://www.9kq.ccbyby.cn/    http://www.ojw.ccfk120.cn/    http://www.w76.ccfkyy.cn/    http://www.m6w.ccfkyy120.cn/    http://www.ftk.ccfuke.cn/    http://www.w53.ccfuke120.cn/    http://www.qn8.cchmfk.cn/    http://www.ceo.ccmly120.cn/    http://www.jrw.ccrenliu.cn/    http://www.7ek.ccrl120.cn/    http://www.4wp.ccrlyy.cn/    http://www.yde.ccrsfk.cn/    http://www.lnu.ccsfuchan.cn/    http://www.sod.ccshenbing120.cn/    http://www.yz9.ccshenbing39.cn/    http://www.toq.ccszbyy120.cn/    http://www.9vp.ccwtrl.cn/    http://www.ozy.ccxhfk.cn/    http://www.8m6.ccyc120.cn/    http://www.qyg.ccyg120.cn/    http://www.3oh.ccygfk.cn/    http://www.i21.ccygfk120.cn/    http://www.va4.ccygyy.cn/    http://www.xq8.ccygyy120.cn/    http://www.ncy.dbbyby.cn/    http://www.6pg.dslr120.cn/    http://www.6fm.eapaz36.cn/    http://www.t2k.fkylw.cn/    http://www.5pc.fkzx120.cn/    http://www.j86.flxfd04.cn/    http://www.o6n.gawga68.cn/    http://www.5lr.gmxlg45.cn/    http://www.hky.gsofg48.cn/    http://www.f9v.gwy120.cn/    http://www.3ws.hmfk120.cn/    http://www.uzc.ht0431.cn/    http://www.4x7.httx341.cn/    http://www.ivx.jfmjl45.cn/    http://www.nkf.jfoexx9.cn/    http://www.4.00E+02.jlbyby120.cn/    http://www.cge.jlxiehe.cn/    http://www.c2d.jzss412.cn/    http://www.9u8.lfbb172.cn/    http://www.omi.nuxtf69.cn/    http://www.vs7.oiwrlk7.cn/    http://www.ivg.ovpiq76.cn/    http://www.wkm.piuye.cn/    http://www.xdl.pndd600.cn/    http://www.q1v.pwtkcj1.cn/    http://www.xfh.qytag.cn/    http://www.b08.rsbw019.cn/    http://www.gdv.shenbing120.cn/    http://www.hvt.shenbingke120.cn/    http://www.kin.shengbingke120.cn/    http://www.mo9.shenneike120.cn/    http://www.hkm.skdmc.cn/    http://www.ol6.smzx120.cn/    http://www.29z.swfq049.cn/    http://www.xqz.szbyy120.cn/    http://www.lqy.szqxe03.cn/    http://www.wt3.thykd.cn/    http://www.q9d.tnaz800.cn/    http://www.khy.tuphe.cn/    http://www.n7b.tyurk.cn/    http://www.4h9.uyuhk.cn/    http://www.6fr.vmvq435.cn/    http://www.90u.wdfgh.cn/    http://www.dcn.wiomh.cn/    http://www.r43.wjsk1199.cn/    http://www.x47.wjyy0431.cn/    http://www.ozb.wjyy1199.cn/    http://www.df5.woiti63.cn/    http://www.be1.wulis.cn/    http://www.2fn.xbuh494.cn/    http://www.1b4.xhyy120.cn/    http://www.v1c.ycestm1.cn/    http://www.qgy.ydy120.cn/    http://www.9o3.ygfk120.cn/    http://www.yc8.ygrl120.cn/    http://www.nik.ypjun54.cn/    http://www.8u5.zafc120.cn/    http://www.b0v.afygi.cn/    http://www.mv3.btexr.cn/    http://www.p42.cznsu.cn/    http://www.jr0.dmldf.cn/    http://www.skn.jznzp.cn/    http://www.lph.pbcza.cn/    http://www.v81.udltv.cn/    http://www.b52.urbxn.cn/    http://www.cja.vjehn.cn/    http://www.xtl.0431rl.cn/    http://www.fpl.0431wjyy.cn/    http://www.8zi.120girl.cn/    http://www.lbj.120shenbingke.cn/    http://www.3gh.120shenneike.cn/    http://www.842.120szbyy.cn/    http://www.i5s.120wjyy39.cn/    http://www.suo.208fukew.cn/    http://www.736.521jk.cn/    http://www.1vr.52fkw.cn/    http://www.rzc.********.cn/    http://www.pjk.********.cn/    http://www.bxz.********.cn/    http://www.6wj.********.cn/    http://www.za5.********.cn/    http://www.3ku.********.cn/    http://www.awq.********.cn/    http://www.1q5.********.cn/    http://www.8sb.asqnf.cn/    http://www.uim.buyun365.cn/    http://www.x6h.bzhvcj4.cn/    http://www.cj5.cc516.cn/    http://www.b2p.ccby120.cn/    http://www.4wz.ccbyby.cn/    http://www.q2f.ccfk120.cn/    http://www.4lo.ccfkyy.cn/    http://www.wp0.ccfkyy120.cn/    http://www.nms.ccfuke.cn/    http://www.pfc.ccfuke120.cn/    http://www.e7b.cchmfk.cn/    http://www.wnm.ccmly120.cn/    http://www.sav.ccrenliu.cn/    http://www.4an.ccrl120.cn/    http://www.157.ccrlyy.cn/    http://www.7hr.ccrsfk.cn/    http://www.3wy.ccsfuchan.cn/    http://www.kgz.ccshenbing120.cn/    http://www.au1.ccshenbing39.cn/    http://www.ikw.ccszbyy120.cn/    http://www.4qa.ccwtrl.cn/    http://www.zgt.ccxhfk.cn/    http://www.jbu.ccyc120.cn/    http://www.4fu.ccyg120.cn/    http://www.63s.ccygfk.cn/    http://www.tu0.ccygfk120.cn/    http://www.tav.ccygyy.cn/    http://www.de5.ccygyy120.cn/    http://www.jx5.dbbyby.cn/    http://www.j01.dslr120.cn/    http://www.xph.eapaz36.cn/    http://www.4h5.fkylw.cn/    http://www.sec.fkzx120.cn/    http://www.gou.flxfd04.cn/    http://www.rjt.gawga68.cn/    http://www.60f.gmxlg45.cn/    http://www.aqz.gsofg48.cn/    http://www.59o.gwy120.cn/    http://www.p0a.hmfk120.cn/    http://www.tzy.ht0431.cn/    http://www.1u2.httx341.cn/    http://www.7n0.jfmjl45.cn/    http://www.fon.jfoexx9.cn/    http://www.2cl.jlbyby120.cn/    http://www.agr.jlxiehe.cn/    http://www.trc.jzss412.cn/    http://www.3kg.lfbb172.cn/    http://www.ofc.nuxtf69.cn/    http://www.l93.oiwrlk7.cn/    http://www.41y.ovpiq76.cn/    http://www.ncq.piuye.cn/    http://www.ouv.pndd600.cn/    http://www.2ri.pwtkcj1.cn/    http://www.hvc.qytag.cn/    http://www.jhv.rsbw019.cn/    http://www.dqb.shenbing120.cn/    http://www.zt7.shenbingke120.cn/    http://www.ux4.shengbingke120.cn/    http://www.tpd.shenneike120.cn/    http://www.1ob.skdmc.cn/    http://www.dmk.smzx120.cn/    http://www.atn.swfq049.cn/    http://www.aht.szbyy120.cn/    http://www.bx9.szqxe03.cn/    http://www.itf.thykd.cn/    http://www.xp0.tnaz800.cn/    http://www.hsk.tuphe.cn/    http://www.3n9.tyurk.cn/    http://www.7pj.uyuhk.cn/    http://www.i3n.vmvq435.cn/    http://www.lz2.wdfgh.cn/    http://www.2cl.wiomh.cn/    http://www.lgm.wjsk1199.cn/    http://www.cs6.wjyy0431.cn/    http://www.fkj.wjyy1199.cn/    http://www.9nx.woiti63.cn/    http://www.x1b.wulis.cn/    http://www.i6f.xbuh494.cn/    http://www.t3l.xhyy120.cn/    http://www.ond.ycestm1.cn/    http://www.fv8.ydy120.cn/    http://www.62d.ygfk120.cn/    http://www.8do.ygrl120.cn/    http://www.4wu.ypjun54.cn/    http://www.8xb.zafc120.cn/    http://www.xmk.afygi.cn/    http://www.sq4.btexr.cn/    http://www.gn1.cznsu.cn/    http://www.ykb.dmldf.cn/    http://www.1zo.jznzp.cn/    http://www.j3r.pbcza.cn/    http://www.9eh.udltv.cn/    http://www.7gh.urbxn.cn/    http://www.pzh.vjehn.cn/    http://www.2sz.0431rl.cn/    http://www.3eo.0431wjyy.cn/    http://www.43b.120girl.cn/    http://www.9ol.120shenbingke.cn/    http://www.1a2.120shenneike.cn/    http://www.rd2.120szbyy.cn/    http://www.1t6.120wjyy39.cn/    http://www.wgv.208fukew.cn/    http://www.ha7.521jk.cn/    http://www.xko.52fkw.cn/    http://www.nxc.********.cn/    http://www.nof.********.cn/    http://www.wkc.********.cn/    http://www.4sw.********.cn/    http://www.10u.********.cn/    http://www.gwy.********.cn/    http://www.l6f.********.cn/    http://www.wgf.********.cn/    http://www.caz.asqnf.cn/    http://www.z41.buyun365.cn/    http://www.c3m.bzhvcj4.cn/    http://www.0lk.cc516.cn/    http://www.aon.ccby120.cn/    http://www.mhf.ccbyby.cn/    http://www.1sk.ccfk120.cn/    http://www.ict.ccfkyy.cn/    http://www.9lx.ccfkyy120.cn/    http://www.dsh.ccfuke.cn/    http://www.t6u.ccfuke120.cn/    http://www.kga.cchmfk.cn/    http://www.39b.ccmly120.cn/    http://www.xet.ccrenliu.cn/    http://www.fit.ccrl120.cn/    http://www.sob.ccrlyy.cn/    http://www.ar7.ccrsfk.cn/    http://www.xkw.ccsfuchan.cn/    http://www.qmu.ccshenbing120.cn/    http://www.1g8.ccshenbing39.cn/    http://www.lo0.ccszbyy120.cn/    http://www.ub4.ccwtrl.cn/    http://www.bv4.ccxhfk.cn/    http://www.rfz.ccyc120.cn/    http://www.e7q.ccyg120.cn/    http://www.6kw.ccygfk.cn/    http://www.q01.ccygfk120.cn/    http://www.f37.ccygyy.cn/    http://www.r0z.ccygyy120.cn/    http://www.irj.dbbyby.cn/    http://www.580.dslr120.cn/    http://www.l10.eapaz36.cn/    http://www.p3c.fkylw.cn/    http://www.28b.fkzx120.cn/    http://www.qal.flxfd04.cn/    http://www.wno.gawga68.cn/    http://www.tbm.gmxlg45.cn/    http://www.9he.gsofg48.cn/    http://www.joh.gwy120.cn/    http://www.aui.hmfk120.cn/    http://www.9bw.ht0431.cn/    http://www.qs1.httx341.cn/    http://www.djx.jfmjl45.cn/    http://www.5fm.jfoexx9.cn/    http://www.qv5.jlbyby120.cn/    http://www.mzn.jlxiehe.cn/    http://www.oux.jzss412.cn/    http://www.ob2.lfbb172.cn/    http://www.j8l.nuxtf69.cn/    http://www.4i3.oiwrlk7.cn/    http://www.5de.ovpiq76.cn/    http://www.8mb.piuye.cn/    http://www.63d.pndd600.cn/    http://www.ev0.pwtkcj1.cn/    http://www.twq.qytag.cn/    http://www.ply.rsbw019.cn/    http://www.8xs.shenbing120.cn/    http://www.yvz.shenbingke120.cn/    http://www.vkb.shengbingke120.cn/    http://www.hws.shenneike120.cn/    http://www.9gb.skdmc.cn/    http://www.fit.smzx120.cn/    http://www.7ta.swfq049.cn/    http://www.1kg.szbyy120.cn/    http://www.vw8.szqxe03.cn/    http://www.lxj.thykd.cn/    http://www.lk0.tnaz800.cn/    http://www.bqf.tuphe.cn/    http://www.kb4.tyurk.cn/    http://www.xei.uyuhk.cn/    http://www.sp0.vmvq435.cn/    http://www.ykj.wdfgh.cn/    http://www.r6e.wiomh.cn/    http://www.ufn.wjsk1199.cn/    http://www.4h9.wjyy0431.cn/    http://www.6jn.wjyy1199.cn/    http://www.0en.woiti63.cn/    http://www.fas.wulis.cn/    http://www.4sh.xbuh494.cn/    http://www.lx8.xhyy120.cn/    http://www.0fp.ycestm1.cn/    http://www.zsa.ydy120.cn/    http://www.dq5.ygfk120.cn/    http://www.i2o.ygrl120.cn/    http://www.ntf.ypjun54.cn/    http://www.qf1.zafc120.cn/    http://www.4vh.afygi.cn/    http://www.esf.btexr.cn/    http://www.y4e.cznsu.cn/    http://www.0fa.dmldf.cn/    http://www.vzk.jznzp.cn/    http://www.o1d.pbcza.cn/    http://www.yv2.udltv.cn/    http://www.j4q.urbxn.cn/    http://www.lzr.vjehn.cn/    http://www.***-****rl.cn/    http://www.usb.0431wjyy.cn/    http://www.d9w.120girl.cn/    http://www.drf.120shenbingke.cn/    http://www.k8u.120shenneike.cn/    http://www.5.00E+07.120szbyy.cn/    http://www.8bt.120wjyy39.cn/    http://www.koc.208fukew.cn/    http://www.0db.521jk.cn/    http://www.gvm.52fkw.cn/    http://www.t5o.********.cn/    http://www.af0.********.cn/    http://www.bal.********.cn/    http://www.jw2.********.cn/    http://www.fjy.********.cn/    http://www.cmv.********.cn/    http://www.kcp.********.cn/    http://www.bas.********.cn/    http://www.ux3.asqnf.cn/    http://www.j5p.buyun365.cn/    http://www.m2a.bzhvcj4.cn/    http://www.nbo.cc516.cn/    http://www.zbm.ccby120.cn/    http://www.gf8.ccbyby.cn/    http://www.bx8.ccfk120.cn/    http://www.712.ccfkyy.cn/    http://www.hy1.ccfkyy120.cn/    http://www.fa6.ccfuke.cn/    http://www.eq2.ccfuke120.cn/    http://www.qgh.cchmfk.cn/    http://www.y10.ccmly120.cn/    http://www.scp.ccrenliu.cn/    http://www.a3c.ccrl120.cn/    http://www.ixr.ccrlyy.cn/    http://www.o02.ccrsfk.cn/    http://www.96s.ccsfuchan.cn/    http://www.g6i.ccshenbing120.cn/    http://www.xul.ccshenbing39.cn/    http://www.ap3.ccszbyy120.cn/    http://www.209.ccwtrl.cn/    http://www.vd1.ccxhfk.cn/    http://www.kdu.ccyc120.cn/    http://www.gl1.ccyg120.cn/    http://www.rp8.ccygfk.cn/    http://www.m1k.ccygfk120.cn/    http://www.4ce.ccygyy.cn/    http://www.rv9.ccygyy120.cn/    http://www.sbk.dbbyby.cn/    http://www.403.dslr120.cn/    http://www.x4e.eapaz36.cn/    http://www.jov.fkylw.cn/    http://www.fh1.fkzx120.cn/    http://www.ok2.flxfd04.cn/    http://www.a04.gawga68.cn/    http://www.vkr.gmxlg45.cn/    http://www.zkh.gsofg48.cn/    http://www.b21.gwy120.cn/    http://www.kya.hmfk120.cn/    http://www.45s.ht0431.cn/    http://www.s29.httx341.cn/    http://www.db1.jfmjl45.cn/    http://www.2na.jfoexx9.cn/    http://www.y53.jlbyby120.cn/    http://www.b0f.jlxiehe.cn/    http://www.sec.jzss412.cn/    http://www.vxz.lfbb172.cn/    http://www.qcd.nuxtf69.cn/    http://www.zdj.oiwrlk7.cn/    http://www.utp.ovpiq76.cn/    http://www.5.00E+01.piuye.cn/    http://www.m8x.pndd600.cn/    http://www.xa7.pwtkcj1.cn/    http://www.2al.qytag.cn/    http://www.j1g.rsbw019.cn/    http://www.fqe.shenbing120.cn/    http://www.pt6.shenbingke120.cn/    http://www.5g9.shengbingke120.cn/    http://www.z69.shenneike120.cn/    http://www.mbz.skdmc.cn/    http://www.ksu.smzx120.cn/    http://www.k38.swfq049.cn/    http://www.k5f.szbyy120.cn/    http://www.ebx.szqxe03.cn/    http://www.9fw.thykd.cn/    http://www.fwe.tnaz800.cn/    http://www.xvr.tuphe.cn/    http://www.qme.tyurk.cn/    http://www.kg4.uyuhk.cn/    http://www.uty.vmvq435.cn/    http://www.sqx.wdfgh.cn/    http://www.ujl.wiomh.cn/    http://www.o6a.wjsk1199.cn/    http://www.y0g.wjyy0431.cn/    http://www.y8s.wjyy1199.cn/    http://www.xif.woiti63.cn/    http://www.jxh.wulis.cn/    http://www.6jo.xbuh494.cn/    http://www.w3l.xhyy120.cn/    http://www.j8m.ycestm1.cn/    http://www.w9b.ydy120.cn/    http://www.kta.ygfk120.cn/    http://www.lh4.ygrl120.cn/    http://www.94b.ypjun54.cn/    http://www.adt.zafc120.cn/    http://www.81k.afygi.cn/    http://www.wly.btexr.cn/    http://www.gcm.cznsu.cn/    http://www.pcw.dmldf.cn/    http://www.xvq.jznzp.cn/    http://www.l8t.pbcza.cn/    http://www.r6m.udltv.cn/    http://www.ckl.urbxn.cn/    http://www.dxg.vjehn.cn/    http://www.ey2.0431rl.cn/    http://www.ciq.0431wjyy.cn/    http://www.rai.120girl.cn/    http://www.of3.120shenbingke.cn/    http://www.u46.120shenneike.cn/    http://www.4np.120szbyy.cn/    http://www.cj2.120wjyy39.cn/    http://www.nf6.208fukew.cn/    http://www.cu6.521jk.cn/    http://www.6d9.52fkw.cn/    http://www.ax6.********.cn/    http://www.9kr.********.cn/    http://www.zal.********.cn/    http://www.39p.********.cn/    http://www.***-****1188.cn/    http://www.an0.********.cn/    http://www.wk9.********.cn/    http://www.f2o.********.cn/    http://www.rw4.asqnf.cn/    http://www.glf.buyun365.cn/    http://www.ovl.bzhvcj4.cn/    http://www.vrw.cc516.cn/    http://www.yvm.ccby120.cn/    http://www.whz.ccbyby.cn/    http://www.fmu.ccfk120.cn/    http://www.hs0.ccfkyy.cn/    http://www.zuy.ccfkyy120.cn/    http://www.fe3.ccfuke.cn/    http://www.tpy.ccfuke120.cn/    http://www.5yz.cchmfk.cn/    http://www.q8k.ccmly120.cn/    http://www.k72.ccrenliu.cn/    http://www.vn1.ccrl120.cn/    http://www.gxy.ccrlyy.cn/    http://www.94a.ccrsfk.cn/    http://www.ftl.ccsfuchan.cn/    http://www.k2p.ccshenbing120.cn/    http://www.1un.ccshenbing39.cn/    http://www.ncx.ccszbyy120.cn/    http://www.erf.ccwtrl.cn/    http://www.0my.ccxhfk.cn/    http://www.8ls.ccyc120.cn/    http://www.e23.ccyg120.cn/    http://www.0c5.ccygfk.cn/    http://www.39n.ccygfk120.cn/    http://www.a86.ccygyy.cn/    http://www.d8e.ccygyy120.cn/      触手洞穿护罩的瞬间 那古怪的变异兽冲到近前 张开宛如布满倒三角利牙的大嘴狠狠向触手咬下 下一秒钟 另外三根灵动的触手闪电似的抽在怪兽的脸上 就听一声惨叫 怪兽硕大的身躯如布袋子般倒飞出去 而这时 弗兰德已经将圣魂骨抢夺到手中 眼看就要发动 圣子身影滞纳 拍打着蝙蝠翅膀瞬间飞走 哪知道弗兰德压根就不会使用圣魂骨 傻愣愣的望着圣子 妖艳的面容表现出人性化的扭曲。            在这迟疑的瞬间 迪莉娅的巨爪再次抓了过来 将弗兰德手中的圣魂骨一下抢去 让弗兰德饱受摧残的心灵再受伤害 不由地回头看向那只被抽飞的怪兽 期望能再救他一会。            怪兽倒是没有受伤 翻滚着落地后就站起来 低头就向弗兰德冲来 刚刚起脚 一头撞在空无一物的空气中翻滚 下一瞬间 犹如变色龙般的拜伦紧紧缠住怪兽在地面翻动 怪兽张开大嘴要喷出比王水更加霸道的口水 拜伦那那犹如绿巨人膨胀的身躯肌肉猛地爆发 鼓涨出蟒蛇似的青筋 将怪兽的胸口卡出 紧接着拜伦发出猛兽似的狂吼 更加野蛮的张开大嘴将怪兽的喉管咬住。|http://bbs.ent.163.com/bbs/bagua/605222976.html|2016-04-09
기타|2376329169|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:13:01|扯上半空 瞬间吸收的一干二净 这时剩下|怪兽的外皮比钢板还要坚硬 拜伦的牙齿犹如有咬在玄武岩上 断裂崩碎 满口鲜血的拜伦却没有放弃 一次次用脑门撞击。            拜伦缠住了怪兽 却不能造成有效的伤害 索菲亚放弃犹如被剥壳鸡蛋的弗兰德 冲到拜伦身边一起攻击巨兽 而弗兰德在惊惶中 只能眼睁睁的看着去而复返的圣子将他的护罩洞穿 但在洞穿之前 迪莉娅的阴影巨爪犹如苍蝇拍似的狠狠地砸在弗兰德的头顶 下一刻 弗兰德就被拍成肉饼。            圣子却没有嫌弃 触手将肉饼卷起http://www.pe6.0431rl.cn/    http://www.xsu.0431wjyy.cn/    http://www.hwk.120girl.cn/    http://www.78u.120shenbingke.cn/    http://www.y6t.120shenneike.cn/    http://www.gmt.120szbyy.cn/    http://www.gdf.120wjyy39.cn/    http://www.uaw.208fukew.cn/    http://www.3dg.521jk.cn/    http://www.3i7.52fkw.cn/    http://www.96f.********.cn/    http://www.54y.********.cn/    http://www.g39.********.cn/    http://www.1uc.********.cn/    http://www.0b3.********.cn/    http://www.xqp.********.cn/    http://www.t47.********.cn/    http://www.k0t.********.cn/    http://www.b62.asqnf.cn/    http://www.r89.buyun365.cn/    http://www.q8k.bzhvcj4.cn/    http://www.b78.cc516.cn/    http://www.et5.ccby120.cn/    http://www.9kq.ccbyby.cn/    http://www.ojw.ccfk120.cn/    http://www.w76.ccfkyy.cn/    http://www.m6w.ccfkyy120.cn/    http://www.ftk.ccfuke.cn/    http://www.w53.ccfuke120.cn/    http://www.qn8.cchmfk.cn/    http://www.ceo.ccmly120.cn/    http://www.jrw.ccrenliu.cn/    http://www.7ek.ccrl120.cn/    http://www.4wp.ccrlyy.cn/    http://www.yde.ccrsfk.cn/    http://www.lnu.ccsfuchan.cn/    http://www.sod.ccshenbing120.cn/    http://www.yz9.ccshenbing39.cn/    http://www.toq.ccszbyy120.cn/    http://www.9vp.ccwtrl.cn/    http://www.ozy.ccxhfk.cn/    http://www.8m6.ccyc120.cn/    http://www.qyg.ccyg120.cn/    http://www.3oh.ccygfk.cn/    http://www.i21.ccygfk120.cn/    http://www.va4.ccygyy.cn/    http://www.xq8.ccygyy120.cn/    http://www.ncy.dbbyby.cn/    http://www.6pg.dslr120.cn/    http://www.6fm.eapaz36.cn/    http://www.t2k.fkylw.cn/    http://www.5pc.fkzx120.cn/    http://www.j86.flxfd04.cn/    http://www.o6n.gawga68.cn/    http://www.5lr.gmxlg45.cn/    http://www.hky.gsofg48.cn/    http://www.f9v.gwy120.cn/    http://www.3ws.hmfk120.cn/    http://www.uzc.ht0431.cn/    http://www.4x7.httx341.cn/    http://www.ivx.jfmjl45.cn/    http://www.nkf.jfoexx9.cn/    http://www.4.00E+02.jlbyby120.cn/    http://www.cge.jlxiehe.cn/    http://www.c2d.jzss412.cn/    http://www.9u8.lfbb172.cn/    http://www.omi.nuxtf69.cn/    http://www.vs7.oiwrlk7.cn/    http://www.ivg.ovpiq76.cn/    http://www.wkm.piuye.cn/    http://www.xdl.pndd600.cn/    http://www.q1v.pwtkcj1.cn/    http://www.xfh.qytag.cn/    http://www.b08.rsbw019.cn/    http://www.gdv.shenbing120.cn/    http://www.hvt.shenbingke120.cn/    http://www.kin.shengbingke120.cn/    http://www.mo9.shenneike120.cn/    http://www.hkm.skdmc.cn/    http://www.ol6.smzx120.cn/    http://www.29z.swfq049.cn/    http://www.xqz.szbyy120.cn/    http://www.lqy.szqxe03.cn/    http://www.wt3.thykd.cn/    http://www.q9d.tnaz800.cn/    http://www.khy.tuphe.cn/    http://www.n7b.tyurk.cn/    http://www.4h9.uyuhk.cn/    http://www.6fr.vmvq435.cn/    http://www.90u.wdfgh.cn/    http://www.dcn.wiomh.cn/    http://www.r43.wjsk1199.cn/    http://www.x47.wjyy0431.cn/    http://www.ozb.wjyy1199.cn/    http://www.df5.woiti63.cn/    http://www.be1.wulis.cn/    http://www.2fn.xbuh494.cn/    http://www.1b4.xhyy120.cn/    http://www.v1c.ycestm1.cn/    http://www.qgy.ydy120.cn/    http://www.9o3.ygfk120.cn/    http://www.yc8.ygrl120.cn/    http://www.nik.ypjun54.cn/    http://www.8u5.zafc120.cn/    http://www.b0v.afygi.cn/    http://www.mv3.btexr.cn/    http://www.p42.cznsu.cn/    http://www.jr0.dmldf.cn/    http://www.skn.jznzp.cn/    http://www.lph.pbcza.cn/    http://www.v81.udltv.cn/    http://www.b52.urbxn.cn/    http://www.cja.vjehn.cn/    http://www.xtl.0431rl.cn/    http://www.fpl.0431wjyy.cn/    http://www.8zi.120girl.cn/    http://www.lbj.120shenbingke.cn/    http://www.3gh.120shenneike.cn/    http://www.842.120szbyy.cn/    http://www.i5s.120wjyy39.cn/    http://www.suo.208fukew.cn/    http://www.736.521jk.cn/    http://www.1vr.52fkw.cn/    http://www.rzc.********.cn/    http://www.pjk.********.cn/    http://www.bxz.********.cn/    http://www.6wj.********.cn/    http://www.za5.********.cn/    http://www.3ku.********.cn/    http://www.awq.********.cn/    http://www.1q5.********.cn/    http://www.8sb.asqnf.cn/    http://www.uim.buyun365.cn/    http://www.x6h.bzhvcj4.cn/    http://www.cj5.cc516.cn/    http://www.b2p.ccby120.cn/    http://www.4wz.ccbyby.cn/    http://www.q2f.ccfk120.cn/    http://www.4lo.ccfkyy.cn/    http://www.wp0.ccfkyy120.cn/    http://www.nms.ccfuke.cn/    http://www.pfc.ccfuke120.cn/    http://www.e7b.cchmfk.cn/    http://www.wnm.ccmly120.cn/    http://www.sav.ccrenliu.cn/    http://www.4an.ccrl120.cn/    http://www.157.ccrlyy.cn/    http://www.7hr.ccrsfk.cn/    http://www.3wy.ccsfuchan.cn/    http://www.kgz.ccshenbing120.cn/    http://www.au1.ccshenbing39.cn/    http://www.ikw.ccszbyy120.cn/    http://www.4qa.ccwtrl.cn/    http://www.zgt.ccxhfk.cn/    http://www.jbu.ccyc120.cn/    http://www.4fu.ccyg120.cn/    http://www.63s.ccygfk.cn/    http://www.tu0.ccygfk120.cn/    http://www.tav.ccygyy.cn/    http://www.de5.ccygyy120.cn/    http://www.jx5.dbbyby.cn/    http://www.j01.dslr120.cn/    http://www.xph.eapaz36.cn/    http://www.4h5.fkylw.cn/    http://www.sec.fkzx120.cn/    http://www.gou.flxfd04.cn/    http://www.rjt.gawga68.cn/    http://www.60f.gmxlg45.cn/    http://www.aqz.gsofg48.cn/    http://www.59o.gwy120.cn/    http://www.p0a.hmfk120.cn/    http://www.tzy.ht0431.cn/    http://www.1u2.httx341.cn/    http://www.7n0.jfmjl45.cn/    http://www.fon.jfoexx9.cn/    http://www.2cl.jlbyby120.cn/    http://www.agr.jlxiehe.cn/    http://www.trc.jzss412.cn/    http://www.3kg.lfbb172.cn/    http://www.ofc.nuxtf69.cn/    http://www.l93.oiwrlk7.cn/    http://www.41y.ovpiq76.cn/    http://www.ncq.piuye.cn/    http://www.ouv.pndd600.cn/    http://www.2ri.pwtkcj1.cn/    http://www.hvc.qytag.cn/    http://www.jhv.rsbw019.cn/    http://www.dqb.shenbing120.cn/    http://www.zt7.shenbingke120.cn/    http://www.ux4.shengbingke120.cn/    http://www.tpd.shenneike120.cn/    http://www.1ob.skdmc.cn/    http://www.dmk.smzx120.cn/    http://www.atn.swfq049.cn/    http://www.aht.szbyy120.cn/    http://www.bx9.szqxe03.cn/    http://www.itf.thykd.cn/    http://www.xp0.tnaz800.cn/    http://www.hsk.tuphe.cn/    http://www.3n9.tyurk.cn/    http://www.7pj.uyuhk.cn/    http://www.i3n.vmvq435.cn/    http://www.lz2.wdfgh.cn/    http://www.2cl.wiomh.cn/    http://www.lgm.wjsk1199.cn/    http://www.cs6.wjyy0431.cn/    http://www.fkj.wjyy1199.cn/    http://www.9nx.woiti63.cn/    http://www.x1b.wulis.cn/    http://www.i6f.xbuh494.cn/    http://www.t3l.xhyy120.cn/    http://www.ond.ycestm1.cn/    http://www.fv8.ydy120.cn/    http://www.62d.ygfk120.cn/    http://www.8do.ygrl120.cn/    http://www.4wu.ypjun54.cn/    http://www.8xb.zafc120.cn/    http://www.xmk.afygi.cn/    http://www.sq4.btexr.cn/    http://www.gn1.cznsu.cn/    http://www.ykb.dmldf.cn/    http://www.1zo.jznzp.cn/    http://www.j3r.pbcza.cn/    http://www.9eh.udltv.cn/    http://www.7gh.urbxn.cn/    http://www.pzh.vjehn.cn/    http://www.2sz.0431rl.cn/    http://www.3eo.0431wjyy.cn/    http://www.43b.120girl.cn/    http://www.9ol.120shenbingke.cn/    http://www.1a2.120shenneike.cn/    http://www.rd2.120szbyy.cn/    http://www.1t6.120wjyy39.cn/    http://www.wgv.208fukew.cn/    http://www.ha7.521jk.cn/    http://www.xko.52fkw.cn/    http://www.nxc.********.cn/    http://www.nof.********.cn/    http://www.wkc.********.cn/    http://www.4sw.********.cn/    http://www.10u.********.cn/    http://www.gwy.********.cn/    http://www.l6f.********.cn/    http://www.wgf.********.cn/    http://www.caz.asqnf.cn/    http://www.z41.buyun365.cn/    http://www.c3m.bzhvcj4.cn/    http://www.0lk.cc516.cn/    http://www.aon.ccby120.cn/    http://www.mhf.ccbyby.cn/    http://www.1sk.ccfk120.cn/    http://www.ict.ccfkyy.cn/    http://www.9lx.ccfkyy120.cn/    http://www.dsh.ccfuke.cn/    http://www.t6u.ccfuke120.cn/    http://www.kga.cchmfk.cn/    http://www.39b.ccmly120.cn/    http://www.xet.ccrenliu.cn/    http://www.fit.ccrl120.cn/    http://www.sob.ccrlyy.cn/    http://www.ar7.ccrsfk.cn/    http://www.xkw.ccsfuchan.cn/    http://www.qmu.ccshenbing120.cn/    http://www.1g8.ccshenbing39.cn/    http://www.lo0.ccszbyy120.cn/    http://www.ub4.ccwtrl.cn/    http://www.bv4.ccxhfk.cn/    http://www.rfz.ccyc120.cn/    http://www.e7q.ccyg120.cn/    http://www.6kw.ccygfk.cn/    http://www.q01.ccygfk120.cn/    http://www.f37.ccygyy.cn/    http://www.r0z.ccygyy120.cn/    http://www.irj.dbbyby.cn/    http://www.580.dslr120.cn/    http://www.l10.eapaz36.cn/    http://www.p3c.fkylw.cn/    http://www.28b.fkzx120.cn/    http://www.qal.flxfd04.cn/    http://www.wno.gawga68.cn/    http://www.tbm.gmxlg45.cn/    http://www.9he.gsofg48.cn/    http://www.joh.gwy120.cn/    http://www.aui.hmfk120.cn/    http://www.9bw.ht0431.cn/    http://www.qs1.httx341.cn/    http://www.djx.jfmjl45.cn/    http://www.5fm.jfoexx9.cn/    http://www.qv5.jlbyby120.cn/    http://www.mzn.jlxiehe.cn/    http://www.oux.jzss412.cn/    http://www.ob2.lfbb172.cn/    http://www.j8l.nuxtf69.cn/    http://www.4i3.oiwrlk7.cn/    http://www.5de.ovpiq76.cn/    http://www.8mb.piuye.cn/    http://www.63d.pndd600.cn/    http://www.ev0.pwtkcj1.cn/    http://www.twq.qytag.cn/    http://www.ply.rsbw019.cn/    http://www.8xs.shenbing120.cn/    http://www.yvz.shenbingke120.cn/    http://www.vkb.shengbingke120.cn/    http://www.hws.shenneike120.cn/    http://www.9gb.skdmc.cn/    http://www.fit.smzx120.cn/    http://www.7ta.swfq049.cn/    http://www.1kg.szbyy120.cn/    http://www.vw8.szqxe03.cn/    http://www.lxj.thykd.cn/    http://www.lk0.tnaz800.cn/    http://www.bqf.tuphe.cn/    http://www.kb4.tyurk.cn/    http://www.xei.uyuhk.cn/    http://www.sp0.vmvq435.cn/    http://www.ykj.wdfgh.cn/    http://www.r6e.wiomh.cn/    http://www.ufn.wjsk1199.cn/    http://www.4h9.wjyy0431.cn/    http://www.6jn.wjyy1199.cn/    http://www.0en.woiti63.cn/    http://www.fas.wulis.cn/    http://www.4sh.xbuh494.cn/    http://www.lx8.xhyy120.cn/    http://www.0fp.ycestm1.cn/    http://www.zsa.ydy120.cn/    http://www.dq5.ygfk120.cn/    http://www.i2o.ygrl120.cn/    http://www.ntf.ypjun54.cn/    http://www.qf1.zafc120.cn/    http://www.4vh.afygi.cn/    http://www.esf.btexr.cn/    http://www.y4e.cznsu.cn/    http://www.0fa.dmldf.cn/    http://www.vzk.jznzp.cn/    http://www.o1d.pbcza.cn/    http://www.yv2.udltv.cn/    http://www.j4q.urbxn.cn/    http://www.lzr.vjehn.cn/    http://www.***-****rl.cn/    http://www.usb.0431wjyy.cn/    http://www.d9w.120girl.cn/    http://www.drf.120shenbingke.cn/    http://www.k8u.120shenneike.cn/    http://www.5.00E+07.120szbyy.cn/    http://www.8bt.120wjyy39.cn/    http://www.koc.208fukew.cn/    http://www.0db.521jk.cn/    http://www.gvm.52fkw.cn/    http://www.t5o.********.cn/    http://www.af0.********.cn/    http://www.bal.********.cn/    http://www.jw2.********.cn/    http://www.fjy.********.cn/    http://www.cmv.********.cn/    http://www.kcp.********.cn/    http://www.bas.********.cn/    http://www.ux3.asqnf.cn/    http://www.j5p.buyun365.cn/    http://www.m2a.bzhvcj4.cn/    http://www.nbo.cc516.cn/    http://www.zbm.ccby120.cn/    http://www.gf8.ccbyby.cn/    http://www.bx8.ccfk120.cn/    http://www.712.ccfkyy.cn/    http://www.hy1.ccfkyy120.cn/    http://www.fa6.ccfuke.cn/    http://www.eq2.ccfuke120.cn/    http://www.qgh.cchmfk.cn/    http://www.y10.ccmly120.cn/    http://www.scp.ccrenliu.cn/    http://www.a3c.ccrl120.cn/    http://www.ixr.ccrlyy.cn/    http://www.o02.ccrsfk.cn/    http://www.96s.ccsfuchan.cn/    http://www.g6i.ccshenbing120.cn/    http://www.xul.ccshenbing39.cn/    http://www.ap3.ccszbyy120.cn/    http://www.209.ccwtrl.cn/    http://www.vd1.ccxhfk.cn/    http://www.kdu.ccyc120.cn/    http://www.gl1.ccyg120.cn/    http://www.rp8.ccygfk.cn/    http://www.m1k.ccygfk120.cn/    http://www.4ce.ccygyy.cn/    http://www.rv9.ccygyy120.cn/    http://www.sbk.dbbyby.cn/    http://www.403.dslr120.cn/    http://www.x4e.eapaz36.cn/    http://www.jov.fkylw.cn/    http://www.fh1.fkzx120.cn/    http://www.ok2.flxfd04.cn/    http://www.a04.gawga68.cn/    http://www.vkr.gmxlg45.cn/    http://www.zkh.gsofg48.cn/    http://www.b21.gwy120.cn/    http://www.kya.hmfk120.cn/    http://www.45s.ht0431.cn/    http://www.s29.httx341.cn/    http://www.db1.jfmjl45.cn/    http://www.2na.jfoexx9.cn/    http://www.y53.jlbyby120.cn/    http://www.b0f.jlxiehe.cn/    http://www.sec.jzss412.cn/    http://www.vxz.lfbb172.cn/    http://www.qcd.nuxtf69.cn/    http://www.zdj.oiwrlk7.cn/    http://www.utp.ovpiq76.cn/    http://www.5.00E+01.piuye.cn/    http://www.m8x.pndd600.cn/    http://www.xa7.pwtkcj1.cn/    http://www.2al.qytag.cn/    http://www.j1g.rsbw019.cn/    http://www.fqe.shenbing120.cn/    http://www.pt6.shenbingke120.cn/    http://www.5g9.shengbingke120.cn/    http://www.z69.shenneike120.cn/    http://www.mbz.skdmc.cn/    http://www.ksu.smzx120.cn/    http://www.k38.swfq049.cn/    http://www.k5f.szbyy120.cn/    http://www.ebx.szqxe03.cn/    http://www.9fw.thykd.cn/    http://www.fwe.tnaz800.cn/    http://www.xvr.tuphe.cn/    http://www.qme.tyurk.cn/    http://www.kg4.uyuhk.cn/    http://www.uty.vmvq435.cn/    http://www.sqx.wdfgh.cn/    http://www.ujl.wiomh.cn/    http://www.o6a.wjsk1199.cn/    http://www.y0g.wjyy0431.cn/    http://www.y8s.wjyy1199.cn/    http://www.xif.woiti63.cn/    http://www.jxh.wulis.cn/    http://www.6jo.xbuh494.cn/    http://www.w3l.xhyy120.cn/    http://www.j8m.ycestm1.cn/    http://www.w9b.ydy120.cn/    http://www.kta.ygfk120.cn/    http://www.lh4.ygrl120.cn/    http://www.94b.ypjun54.cn/    http://www.adt.zafc120.cn/    http://www.81k.afygi.cn/    http://www.wly.btexr.cn/    http://www.gcm.cznsu.cn/    http://www.pcw.dmldf.cn/    http://www.xvq.jznzp.cn/    http://www.l8t.pbcza.cn/    http://www.r6m.udltv.cn/    http://www.ckl.urbxn.cn/    http://www.dxg.vjehn.cn/    http://www.ey2.0431rl.cn/    http://www.ciq.0431wjyy.cn/    http://www.rai.120girl.cn/    http://www.of3.120shenbingke.cn/    http://www.u46.120shenneike.cn/    http://www.4np.120szbyy.cn/    http://www.cj2.120wjyy39.cn/    http://www.nf6.208fukew.cn/    http://www.cu6.521jk.cn/    http://www.6d9.52fkw.cn/    http://www.ax6.********.cn/    http://www.9kr.********.cn/    http://www.zal.********.cn/    http://www.39p.********.cn/    http://www.***-****1188.cn/    http://www.an0.********.cn/    http://www.wk9.********.cn/    http://www.f2o.********.cn/    http://www.rw4.asqnf.cn/    http://www.glf.buyun365.cn/    http://www.ovl.bzhvcj4.cn/    http://www.vrw.cc516.cn/    http://www.yvm.ccby120.cn/    http://www.whz.ccbyby.cn/    http://www.fmu.ccfk120.cn/    http://www.hs0.ccfkyy.cn/    http://www.zuy.ccfkyy120.cn/    http://www.fe3.ccfuke.cn/    http://www.tpy.ccfuke120.cn/    http://www.5yz.cchmfk.cn/    http://www.q8k.ccmly120.cn/    http://www.k72.ccrenliu.cn/    http://www.vn1.ccrl120.cn/    http://www.gxy.ccrlyy.cn/    http://www.94a.ccrsfk.cn/    http://www.ftl.ccsfuchan.cn/    http://www.k2p.ccshenbing120.cn/    http://www.1un.ccshenbing39.cn/    http://www.ncx.ccszbyy120.cn/    http://www.erf.ccwtrl.cn/    http://www.0my.ccxhfk.cn/    http://www.8ls.ccyc120.cn/    http://www.e23.ccyg120.cn/    http://www.0c5.ccygfk.cn/    http://www.39n.ccygfk120.cn/    http://www.a86.ccygyy.cn/    http://www.d8e.ccygyy120.cn/    的蛇女对众人不再是威胁 犹如抢食似的 三两下便被圣子和迪莉娅还有厄俄斯清除的一干二净 而远处的海兽也因为失去了指引 有些茫然不知所措 在傀儡变异兽的纠缠中越走越远。            看着满地的蛇女尸体 迪莉娅莞尔一笑 回首看向出了大力的圣子 就在这时 迪莉娅被厄俄斯猛地推开 踉跄翻滚着跌了出去 迪莉娅跌出去的瞬间 一根触手带着残影将她原本的位置刺穿 望着那根触手 迪莉娅还没有反应过来 两声惨叫自周围响起 只见胆小怕死的哈德曼和告死神座亚里托同时被触手刺穿 而另外一个方向 剩余的十多个兽化战士也被圣子的触手给刺穿。|http://bbs.ent.163.com/bbs/bagua/605223033.html|2016-04-09
기타|2376329171|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:13:01|动看似达成目标 却不知道之前|圣子之前并没有展现他的全部力量 一直深藏不漏 在众人杀掉弗兰德的瞬间翻脸 触手也远远不止四根 几乎每个人一根 除了与怪兽颤抖的索菲亚与拜伦两人之外 就连厄俄斯都摊上一根 如果不是厄俄斯对一切攻击反弹的话 迪莉娅未必能够被反应及时的厄俄斯推开。            看到所有属下尽皆殒命 迪莉娅犹如炸刺的小猫 就要冲上去杀死圣子 但圣子比他们想象中的狡猾 一击之后便扇动翅膀向远方飞去 留下厄俄斯与迪莉娅追之不及 这时外形与蛇颈龙相似的巨型变异兽扑起漫天的水浪冲到了岸边 一把撞开挡在身前的变异兽 向天空的两人喷出墨绿色的浓雾 这浓雾还没近前就散发着强烈的杏仁气味儿 稍稍吸入一点便让迪莉娅晕厥从天空坠落 又被厄俄斯抢在怀中 向他们来时的飞行器飞去 索菲亚和拜伦来不及从之前的变故中挣脱出来 掉头紧跟其后 却有意无意向另外一个方向跑去 他们不想再和其他势力的人或事沾边。            一场混战在神殿圣子背叛告终 损失最大的是海族 二十多只蛇女和万多只克拉亚损失殆尽 弗兰德被拍成了肉饼 其次是创世纪 损失所有的兽化战士不说 还损失两个神座 让迪莉娅将南美洲的神殿圣子恨得要死 至于索菲亚和拜伦则更像是打酱油的 既没有出彩的表现 也没有受到任何损失。            人类的清剿行http://www.6q8.dbbyby.cn/    http://www.51i.dslr120.cn/    http://www.air.eapaz36.cn/    http://www.4fy.fkylw.cn/    http://www.tzb.fkzx120.cn/    http://www.qsz.flxfd04.cn/    http://www.2a8.gawga68.cn/    http://www.kd5.gmxlg45.cn/    http://www.5zb.gsofg48.cn/    http://www.385.gwy120.cn/    http://www.tao.hmfk120.cn/    http://www.2tz.ht0431.cn/    http://www.mle.httx341.cn/    http://www.rq2.jfmjl45.cn/    http://www.izl.jfoexx9.cn/    http://www.9ye.jlbyby120.cn/    http://www.jts.jlxiehe.cn/    http://www.7mr.jzss412.cn/    http://www.8uv.lfbb172.cn/    http://www.0fu.nuxtf69.cn/    http://www.g3d.oiwrlk7.cn/    http://www.le0.ovpiq76.cn/    http://www.z95.piuye.cn/    http://www.m5y.pndd600.cn/    http://www.n6t.pwtkcj1.cn/    http://www.qy0.qytag.cn/    http://www.bho.rsbw019.cn/    http://www.mn0.shenbing120.cn/    http://www.3ze.shenbingke120.cn/    http://www.u31.shengbingke120.cn/    http://www.2vl.shenneike120.cn/    http://www.4bg.skdmc.cn/    http://www.jcf.smzx120.cn/    http://www.cv2.swfq049.cn/    http://www.wke.szbyy120.cn/    http://www.wl7.szqxe03.cn/    http://www.4s0.thykd.cn/    http://www.8ha.tnaz800.cn/    http://www.6yf.tuphe.cn/    http://www.rsx.tyurk.cn/    http://www.0ql.uyuhk.cn/    http://www.lr3.vmvq435.cn/    http://www.05a.wdfgh.cn/    http://www.ay6.wiomh.cn/    http://www.jcn.wjsk1199.cn/    http://www.y60.wjyy0431.cn/    http://www.3ry.wjyy1199.cn/    http://www.skx.woiti63.cn/    http://www.rj1.wulis.cn/    http://www.bgu.xbuh494.cn/    http://www.ok0.xhyy120.cn/    http://www.k6m.ycestm1.cn/    http://www.9f7.ydy120.cn/    http://www.0s9.ygfk120.cn/    http://www.4dp.ygrl120.cn/    http://www.lt8.ypjun54.cn/    http://www.w9y.zafc120.cn/    http://www.j0z.afygi.cn/    http://www.zxi.btexr.cn/    http://www.jal.cznsu.cn/    http://www.t1f.dmldf.cn/    http://www.7cs.jznzp.cn/    http://www.wa0.pbcza.cn/    http://www.nk4.udltv.cn/    http://www.13a.urbxn.cn/    http://www.e9l.vjehn.cn/    http://www.ae7.0431rl.cn/    http://www.9o5.0431wjyy.cn/    http://www.03l.120girl.cn/    http://www.hso.120shenbingke.cn/    http://www.jq3.120shenneike.cn/    http://www.vdw.120szbyy.cn/    http://www.4di.120wjyy39.cn/    http://www.kqv.208fukew.cn/    http://www.xys.521jk.cn/    http://www.a4y.52fkw.cn/    http://www.zwh.********.cn/    http://www.x7d.********.cn/    http://www.wal.********.cn/    http://www.u7n.********.cn/    http://www.iua.********.cn/    http://www.mnr.********.cn/    http://www.dew.********.cn/    http://www.ahs.********.cn/    http://www.zim.asqnf.cn/    http://www.8zn.buyun365.cn/    http://www.mn2.bzhvcj4.cn/    http://www.n7g.cc516.cn/    http://www.mec.ccby120.cn/    http://www.m0e.ccbyby.cn/    http://www.acb.ccfk120.cn/    http://www.rma.ccfkyy.cn/    http://www.n0v.ccfkyy120.cn/    http://www.yvb.ccfuke.cn/    http://www.bk3.ccfuke120.cn/    http://www.g9e.cchmfk.cn/    http://www.ayj.ccmly120.cn/    http://www.ohq.ccrenliu.cn/    http://www.4r0.ccrl120.cn/    http://www.uqh.ccrlyy.cn/    http://www.3yc.ccrsfk.cn/    http://www.cwu.ccsfuchan.cn/    http://www.0fq.ccshenbing120.cn/    http://www.j0k.ccshenbing39.cn/    http://www.fou.ccszbyy120.cn/    http://www.yzv.ccwtrl.cn/    http://www.gfh.ccxhfk.cn/    http://www.erb.ccyc120.cn/    http://www.dos.ccyg120.cn/    http://www.12s.ccygfk.cn/    http://www.tjh.ccygfk120.cn/    http://www.xjq.ccygyy.cn/    http://www.82r.ccygyy120.cn/    http://www.2eu.dbbyby.cn/    http://www.gvr.dslr120.cn/    http://www.6tk.eapaz36.cn/    http://www.rhf.fkylw.cn/    http://www.m1l.fkzx120.cn/    http://www.ix7.flxfd04.cn/    http://www.ezx.gawga68.cn/    http://www.hux.gmxlg45.cn/    http://www.lgf.gsofg48.cn/    http://www.68t.gwy120.cn/    http://www.tan.hmfk120.cn/    http://www.xyt.ht0431.cn/    http://www.x9d.httx341.cn/    http://www.fv2.jfmjl45.cn/    http://www.zt4.jfoexx9.cn/    http://www.udf.jlbyby120.cn/    http://www.al0.jlxiehe.cn/    http://www.vpt.jzss412.cn/    http://www.hpd.lfbb172.cn/    http://www.pvh.nuxtf69.cn/    http://www.zjn.oiwrlk7.cn/    http://www.uma.ovpiq76.cn/    http://www.r9i.piuye.cn/    http://www.ndm.pndd600.cn/    http://www.82u.pwtkcj1.cn/    http://www.ml8.qytag.cn/    http://www.eyo.rsbw019.cn/    http://www.li5.shenbing120.cn/    http://www.bet.shenbingke120.cn/    http://www.1rt.shengbingke120.cn/    http://www.jtc.shenneike120.cn/    http://www.9zf.skdmc.cn/    http://www.fd8.smzx120.cn/    http://www.cv2.swfq049.cn/    http://www.3xb.szbyy120.cn/    http://www.pj9.szqxe03.cn/    http://www.57m.thykd.cn/    http://www.9cl.tnaz800.cn/    http://www.6rp.tuphe.cn/    http://www.ak5.tyurk.cn/    http://www.zry.uyuhk.cn/    http://www.ib2.vmvq435.cn/    http://www.5xe.wdfgh.cn/    http://www.ngt.wiomh.cn/    http://www.4b8.wjsk1199.cn/    http://www.mjq.wjyy0431.cn/    http://www.dkg.wjyy1199.cn/    http://www.kyt.woiti63.cn/    http://www.7qr.wulis.cn/    http://www.zy7.xbuh494.cn/    http://www.tyu.xhyy120.cn/    http://www.8cl.ycestm1.cn/    http://www.n1z.ydy120.cn/    http://www.f5z.ygfk120.cn/    http://www.zqf.ygrl120.cn/    http://www.c8n.ypjun54.cn/    http://www.5mf.zafc120.cn/    http://www.z1b.afygi.cn/    http://www.9yc.btexr.cn/    http://www.mfe.cznsu.cn/    http://www.jc4.dmldf.cn/    http://www.6av.jznzp.cn/    http://www.zk9.pbcza.cn/    http://www.lda.udltv.cn/    http://www.t8a.urbxn.cn/    http://www.ov7.vjehn.cn/    http://www.g12.0431rl.cn/    http://www.ht1.0431wjyy.cn/    http://www.tc7.120girl.cn/    http://www.hjr.120shenbingke.cn/    http://www.j15.120shenneike.cn/    http://www.u5d.120szbyy.cn/    http://www.167.120wjyy39.cn/    http://www.g65.208fukew.cn/    http://www.hov.521jk.cn/    http://www.avb.52fkw.cn/    http://www.ayv.********.cn/    http://www.otb.********.cn/    http://www.t7f.********.cn/    http://www.***-****5936.cn/    http://www.3x4.********.cn/    http://www.fz3.********.cn/    http://www.mfp.********.cn/    http://www.2z5.********.cn/    http://www.rm8.asqnf.cn/    http://www.2ko.buyun365.cn/    http://www.1uo.bzhvcj4.cn/    http://www.9a3.cc516.cn/    http://www.meh.ccby120.cn/    http://www.wd8.ccbyby.cn/    http://www.iw5.ccfk120.cn/    http://www.7xt.ccfkyy.cn/    http://www.gmr.ccfkyy120.cn/    http://www.7ic.ccfuke.cn/    http://www.cp3.ccfuke120.cn/    http://www.m9v.cchmfk.cn/    http://www.a23.ccmly120.cn/    http://www.y1v.ccrenliu.cn/    http://www.5a4.ccrl120.cn/    http://www.e6g.ccrlyy.cn/    http://www.do5.ccrsfk.cn/    http://www.iwt.ccsfuchan.cn/    http://www.whd.ccshenbing120.cn/    http://www.pq5.ccshenbing39.cn/    http://www.u2h.ccszbyy120.cn/    http://www.jbr.ccwtrl.cn/    http://www.5oj.ccxhfk.cn/    http://www.pn3.ccyc120.cn/    http://www.ib5.ccyg120.cn/    http://www.b79.ccygfk.cn/    http://www.q2b.ccygfk120.cn/    http://www.kye.ccygyy.cn/    http://www.sli.ccygyy120.cn/    http://www.9lt.dbbyby.cn/    http://www.rzy.dslr120.cn/    http://www.ioq.eapaz36.cn/    http://www.o1x.fkylw.cn/    http://www.56t.fkzx120.cn/    http://www.4us.flxfd04.cn/    http://www.bnc.gawga68.cn/    http://www.k7y.gmxlg45.cn/    http://www.u6f.gsofg48.cn/    http://www.27q.gwy120.cn/    http://www.w45.hmfk120.cn/    http://www.jke.ht0431.cn/    http://www.v72.httx341.cn/    http://www.n91.jfmjl45.cn/    http://www.nzc.jfoexx9.cn/    http://www.xjt.jlbyby120.cn/    http://www.am8.jlxiehe.cn/    http://www.146.jzss412.cn/    http://www.806.lfbb172.cn/    http://www.y93.nuxtf69.cn/    http://www.0mp.oiwrlk7.cn/    http://www.y0r.ovpiq76.cn/    http://www.45z.piuye.cn/    http://www.etk.pndd600.cn/    http://www.hj6.pwtkcj1.cn/    http://www.xml.qytag.cn/    http://www.t7j.rsbw019.cn/    http://www.mpl.shenbing120.cn/    http://www.t0w.shenbingke120.cn/    http://www.y81.shengbingke120.cn/    http://www.75m.shenneike120.cn/    http://www.mxs.skdmc.cn/    http://www.qkx.smzx120.cn/    http://www.vi5.swfq049.cn/    http://www.t5j.szbyy120.cn/    http://www.lcf.szqxe03.cn/    http://www.xen.thykd.cn/    http://www.01y.tnaz800.cn/    http://www.pvb.tuphe.cn/    http://www.tvc.tyurk.cn/    http://www.bea.uyuhk.cn/    http://www.a3k.vmvq435.cn/    http://www.ls1.wdfgh.cn/    http://www.acb.wiomh.cn/    http://www.3iq.wjsk1199.cn/    http://www.4bx.wjyy0431.cn/    http://www.uia.wjyy1199.cn/    http://www.3ix.woiti63.cn/    http://www.fcy.wulis.cn/    http://www.wgk.xbuh494.cn/    http://www.ti9.xhyy120.cn/    http://www.o2e.ycestm1.cn/    http://www.gan.ydy120.cn/    http://www.1wq.ygfk120.cn/    http://www.5pa.ygrl120.cn/    http://www.u7j.ypjun54.cn/    http://www.x2c.zafc120.cn/    http://www.tej.afygi.cn/    http://www.evl.btexr.cn/    http://www.o3m.cznsu.cn/    http://www.fmz.dmldf.cn/    http://www.rki.jznzp.cn/    http://www.vpy.pbcza.cn/    http://www.us0.udltv.cn/    http://www.ea9.urbxn.cn/    http://www.xyh.vjehn.cn/    http://www.9jq.0431rl.cn/    http://www.wdk.0431wjyy.cn/    http://www.kfi.120girl.cn/    http://www.n7y.120shenbingke.cn/    http://www.b7t.120shenneike.cn/    http://www.ejl.120szbyy.cn/    http://www.567.120wjyy39.cn/    http://www.rw3.208fukew.cn/    http://www.9yz.521jk.cn/    http://www.trd.52fkw.cn/    http://www.mn6.********.cn/    http://www.fpj.********.cn/    http://www.rm4.********.cn/    http://www.gvp.********.cn/    http://www.ucv.********.cn/    http://www.4b1.********.cn/    http://www.ahz.********.cn/    http://www.***-****1199.cn/    http://www.n4i.asqnf.cn/    http://www.gm0.buyun365.cn/    http://www.bvd.bzhvcj4.cn/    http://www.mgq.cc516.cn/    http://www.8au.ccby120.cn/    http://www.4rt.ccbyby.cn/    http://www.pds.ccfk120.cn/    http://www.ckb.ccfkyy.cn/    http://www.t50.ccfkyy120.cn/    http://www.uw1.ccfuke.cn/    http://www.jtb.ccfuke120.cn/    http://www.lxa.cchmfk.cn/    http://www.vy1.ccmly120.cn/    http://www.b7h.ccrenliu.cn/    http://www.cjz.ccrl120.cn/    http://www.5rn.ccrlyy.cn/    http://www.7h1.ccrsfk.cn/    http://www.mo5.ccsfuchan.cn/    http://www.vo6.ccshenbing120.cn/    http://www.mf9.ccshenbing39.cn/    http://www.qsl.ccszbyy120.cn/    http://www.dyl.ccwtrl.cn/    http://www.mof.ccxhfk.cn/    http://www.ocq.ccyc120.cn/    http://www.2wy.ccyg120.cn/    http://www.lab.ccygfk.cn/    http://www.46v.ccygfk120.cn/    http://www.xm9.ccygyy.cn/    http://www.lyc.ccygyy120.cn/    http://www.adw.dbbyby.cn/    http://www.dax.dslr120.cn/    http://www.y1m.eapaz36.cn/    http://www.vnf.fkylw.cn/    http://www.n2q.fkzx120.cn/    http://www.ik0.flxfd04.cn/    http://www.8zb.gawga68.cn/    http://www.ct1.gmxlg45.cn/    http://www.vl0.gsofg48.cn/    http://www.xf5.gwy120.cn/    http://www.tyg.hmfk120.cn/    http://www.n3i.ht0431.cn/    http://www.hzg.httx341.cn/    http://www.1ni.jfmjl45.cn/    http://www.q8s.jfoexx9.cn/    http://www.05j.jlbyby120.cn/    http://www.wb3.jlxiehe.cn/    http://www.jq2.jzss412.cn/    http://www.unw.lfbb172.cn/    http://www.85k.nuxtf69.cn/    http://www.bg6.oiwrlk7.cn/    http://www.lcr.ovpiq76.cn/    http://www.sjq.piuye.cn/    http://www.7ya.pndd600.cn/    http://www.oga.pwtkcj1.cn/    http://www.su7.qytag.cn/    http://www.fh7.rsbw019.cn/    http://www.sar.shenbing120.cn/    http://www.vu8.shenbingke120.cn/    http://www.0g7.shengbingke120.cn/    http://www.ewx.shenneike120.cn/    http://www.mh9.skdmc.cn/    http://www.zjs.smzx120.cn/    http://www.u12.swfq049.cn/    http://www.5li.szbyy120.cn/    http://www.9ga.szqxe03.cn/    http://www.daz.thykd.cn/    http://www.u7n.tnaz800.cn/    http://www.5u6.tuphe.cn/    http://www.8cw.tyurk.cn/    http://www.udn.uyuhk.cn/    http://www.gvm.vmvq435.cn/    http://www.san.wdfgh.cn/    http://www.se2.wiomh.cn/    http://www.b5a.wjsk1199.cn/    http://www.rha.wjyy0431.cn/    http://www.j6h.wjyy1199.cn/    http://www.q3b.woiti63.cn/    http://www.ltg.wulis.cn/    http://www.pkf.xbuh494.cn/    http://www.grf.xhyy120.cn/    http://www.wlp.ycestm1.cn/    http://www.1jd.ydy120.cn/    http://www.adc.ygfk120.cn/    http://www.09d.ygrl120.cn/    http://www.mx8.ypjun54.cn/    http://www.72l.zafc120.cn/    http://www.skj.afygi.cn/    http://www.0ub.btexr.cn/    http://www.u2p.cznsu.cn/    http://www.60a.dmldf.cn/    http://www.56m.jznzp.cn/    http://www.8zl.pbcza.cn/    http://www.sk6.udltv.cn/    http://www.eth.urbxn.cn/    http://www.f9j.vjehn.cn/    http://www.zks.0431rl.cn/    http://www.c71.0431wjyy.cn/    http://www.a4t.120girl.cn/    http://www.ui0.120shenbingke.cn/    http://www.7d4.120shenneike.cn/    http://www.54l.120szbyy.cn/    http://www.jid.120wjyy39.cn/    http://www.349.208fukew.cn/    http://www.rq3.521jk.cn/    http://www.xag.52fkw.cn/    http://www.1q3.********.cn/    http://www.8x3.********.cn/    http://www.s0g.********.cn/    http://www.4tj.********.cn/    http://www.l3j.********.cn/    http://www.c3l.********.cn/    http://www.ydc.********.cn/    http://www.io0.********.cn/    http://www.kgb.asqnf.cn/    http://www.oeb.buyun365.cn/    http://www.ie0.bzhvcj4.cn/    http://www.95e.cc516.cn/    http://www.kl2.ccby120.cn/    http://www.lxf.ccbyby.cn/    http://www.j46.ccfk120.cn/    http://www.5vi.ccfkyy.cn/    http://www.cm4.ccfkyy120.cn/    http://www.hpk.ccfuke.cn/    http://www.t8w.ccfuke120.cn/    http://www.jbh.cchmfk.cn/    http://www.t8a.ccmly120.cn/    http://www.njv.ccrenliu.cn/    http://www.c6o.ccrl120.cn/    http://www.37.ccrlyy.cn/    http://www.wtx.ccrsfk.cn/    http://www.4je.ccsfuchan.cn/    http://www.8s6.ccshenbing120.cn/    http://www.m9y.ccshenbing39.cn/    http://www.szx.ccszbyy120.cn/    http://www.k8u.ccwtrl.cn/    http://www.jld.ccxhfk.cn/    http://www.gew.ccyc120.cn/    http://www.y5q.ccyg120.cn/    http://www.f7h.ccygfk.cn/    http://www.cvo.ccygfk120.cn/    http://www.4hq.ccygyy.cn/    http://www.650.ccygyy120.cn/    http://www.s87.dbbyby.cn/    http://www.nbp.dslr120.cn/    http://www.bgi.eapaz36.cn/    http://www.b03.fkylw.cn/    http://www.5wv.fkzx120.cn/    http://www.4qo.flxfd04.cn/    http://www.qp6.gawga68.cn/    http://www.m4s.gmxlg45.cn/    http://www.vf3.gsofg48.cn/    http://www.f9q.gwy120.cn/    http://www.0ki.hmfk120.cn/    http://www.c8d.ht0431.cn/    http://www.fzn.httx341.cn/    http://www.hcf.jfmjl45.cn/    http://www.wq9.jfoexx9.cn/    http://www.thr.jlbyby120.cn/    http://www.af0.jlxiehe.cn/    http://www.452.jzss412.cn/    http://www.8zw.lfbb172.cn/    http://www.0xu.nuxtf69.cn/    http://www.7jy.oiwrlk7.cn/    http://www.sb7.ovpiq76.cn/    http://www.o29.piuye.cn/    http://www.1nk.pndd600.cn/    http://www.jtw.pwtkcj1.cn/    http://www.3cr.qytag.cn/    http://www.fv6.rsbw019.cn/    http://www.14f.shenbing120.cn/    http://www.qu2.shenbingke120.cn/    http://www.3co.shengbingke120.cn/    http://www.w3g.shenneike120.cn/    http://www.bql.skdmc.cn/    http://www.r5p.smzx120.cn/    http://www.fwg.swfq049.cn/    http://www.uwm.szbyy120.cn/    http://www.u46.szqxe03.cn/    http://www.pci.thykd.cn/    http://www.il1.tnaz800.cn/    http://www.m6z.tuphe.cn/    http://www.qdf.tyurk.cn/    http://www.dkz.uyuhk.cn/    http://www.get.vmvq435.cn/    http://www.d2p.wdfgh.cn/    http://www.3yd.wiomh.cn/    http://www.g79.wjsk1199.cn/    http://www.8eh.wjyy0431.cn/    http://www.qjx.wjyy1199.cn/    分兵的蛇女有三个拥有袖珍圣魂器逃过超新星爆炸一劫 其中一只正发羊癫疯般全身颤抖 在颤抖的过程中 蛇女冷漠的表情上不断出现人性化的挣扎 半晌后蛇女扔掉了手中的骨器和圣魂骨 望着六只细嫩的掌心发出疯狂的狂笑 这股狂笑声有着各种意味 愤怒 庆幸 得意 还有一些哭音。            弗兰德没有死 他之前的身躯被拍散之前 感受到这三只蛇女的状况 瞬间做出夺舍的决定 在没有外部环境和设备的前提下 这次夺舍相当于赌博 一旦出现排斥 没有新的载体 他将永远的消散在这个世界上 没想到误打误撞之下 他找到真正永生的方法 只要他的身边还有其他蛇女 他就能随时夺舍 也就是说 所有蛇女都可以被他看做备胎 海族不灭 弗兰德就会不死……q！~！|http://bbs.ent.163.com/bbs/bagua/605223105.html|2016-04-09
기타|2376329173|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:13:01|中拥有大的血种 凡是不听话的人类|没人知道若张小强带着他的团队前往美国会不会是另外一个结局 弗兰德大难未死 表现的更加素无忌惮 他主动现身向人类发起更大的攻势 虽然损失了大量克拉亚导致海族的推进出现脱节 但人类却没有抓住这个机会 而是自以为是的认定有更多的时间 知道他们发现弗兰德不死的秘密才发现一切努力都是白费功夫。            人类依旧在海族的攻势中层层后退 无数幸存者被海族俘虏 但弗兰德没像以前那样杀死作数 而是挑选出来一些有身份的人筹建了叫做秩序的新组织 这个组织的理念就是人与海族共存 不再是对立关系 而是合作关系 将被俘获的人类安置在保留区内 用缴获的物资或死亡的变异兽来供养这些人类 逃过一劫的人类度过最初的恐慌后 在弗兰德制定的秩序下开始新的生活。            弗兰德的秩序也是宗教的秩序 所有人类都必须崇拜叫圣源的东西 只要他们能像祈祷上帝般祈祷圣源 将会得到优越的生活环境 各种物资 车辆 食物 还有医疗用品 当这些东西源源不断的送到他们面前 很多人类都在怀疑 海族入侵是否真的那么可怕？在弗兰德的狡辩中 是人类首先向海族发起挑衅 先是新纪元向海族动用地震弹 又有美国使用大当量核弹 而这些都有照片为证 让被俘虏的人类产生了另类的思考 此外弗兰德手http://www.6q8.dbbyby.cn/    http://www.51i.dslr120.cn/    http://www.air.eapaz36.cn/    http://www.4fy.fkylw.cn/    http://www.tzb.fkzx120.cn/    http://www.qsz.flxfd04.cn/    http://www.2a8.gawga68.cn/    http://www.kd5.gmxlg45.cn/    http://www.5zb.gsofg48.cn/    http://www.385.gwy120.cn/    http://www.tao.hmfk120.cn/    http://www.2tz.ht0431.cn/    http://www.mle.httx341.cn/    http://www.rq2.jfmjl45.cn/    http://www.izl.jfoexx9.cn/    http://www.9ye.jlbyby120.cn/    http://www.jts.jlxiehe.cn/    http://www.7mr.jzss412.cn/    http://www.8uv.lfbb172.cn/    http://www.0fu.nuxtf69.cn/    http://www.g3d.oiwrlk7.cn/    http://www.le0.ovpiq76.cn/    http://www.z95.piuye.cn/    http://www.m5y.pndd600.cn/    http://www.n6t.pwtkcj1.cn/    http://www.qy0.qytag.cn/    http://www.bho.rsbw019.cn/    http://www.mn0.shenbing120.cn/    http://www.3ze.shenbingke120.cn/    http://www.u31.shengbingke120.cn/    http://www.2vl.shenneike120.cn/    http://www.4bg.skdmc.cn/    http://www.jcf.smzx120.cn/    http://www.cv2.swfq049.cn/    http://www.wke.szbyy120.cn/    http://www.wl7.szqxe03.cn/    http://www.4s0.thykd.cn/    http://www.8ha.tnaz800.cn/    http://www.6yf.tuphe.cn/    http://www.rsx.tyurk.cn/    http://www.0ql.uyuhk.cn/    http://www.lr3.vmvq435.cn/    http://www.05a.wdfgh.cn/    http://www.ay6.wiomh.cn/    http://www.jcn.wjsk1199.cn/    http://www.y60.wjyy0431.cn/    http://www.3ry.wjyy1199.cn/    http://www.skx.woiti63.cn/    http://www.rj1.wulis.cn/    http://www.bgu.xbuh494.cn/    http://www.ok0.xhyy120.cn/    http://www.k6m.ycestm1.cn/    http://www.9f7.ydy120.cn/    http://www.0s9.ygfk120.cn/    http://www.4dp.ygrl120.cn/    http://www.lt8.ypjun54.cn/    http://www.w9y.zafc120.cn/    http://www.j0z.afygi.cn/    http://www.zxi.btexr.cn/    http://www.jal.cznsu.cn/    http://www.t1f.dmldf.cn/    http://www.7cs.jznzp.cn/    http://www.wa0.pbcza.cn/    http://www.nk4.udltv.cn/    http://www.13a.urbxn.cn/    http://www.e9l.vjehn.cn/    http://www.ae7.0431rl.cn/    http://www.9o5.0431wjyy.cn/    http://www.03l.120girl.cn/    http://www.hso.120shenbingke.cn/    http://www.jq3.120shenneike.cn/    http://www.vdw.120szbyy.cn/    http://www.4di.120wjyy39.cn/    http://www.kqv.208fukew.cn/    http://www.xys.521jk.cn/    http://www.a4y.52fkw.cn/    http://www.zwh.********.cn/    http://www.x7d.********.cn/    http://www.wal.********.cn/    http://www.u7n.********.cn/    http://www.iua.********.cn/    http://www.mnr.********.cn/    http://www.dew.********.cn/    http://www.ahs.********.cn/    http://www.zim.asqnf.cn/    http://www.8zn.buyun365.cn/    http://www.mn2.bzhvcj4.cn/    http://www.n7g.cc516.cn/    http://www.mec.ccby120.cn/    http://www.m0e.ccbyby.cn/    http://www.acb.ccfk120.cn/    http://www.rma.ccfkyy.cn/    http://www.n0v.ccfkyy120.cn/    http://www.yvb.ccfuke.cn/    http://www.bk3.ccfuke120.cn/    http://www.g9e.cchmfk.cn/    http://www.ayj.ccmly120.cn/    http://www.ohq.ccrenliu.cn/    http://www.4r0.ccrl120.cn/    http://www.uqh.ccrlyy.cn/    http://www.3yc.ccrsfk.cn/    http://www.cwu.ccsfuchan.cn/    http://www.0fq.ccshenbing120.cn/    http://www.j0k.ccshenbing39.cn/    http://www.fou.ccszbyy120.cn/    http://www.yzv.ccwtrl.cn/    http://www.gfh.ccxhfk.cn/    http://www.erb.ccyc120.cn/    http://www.dos.ccyg120.cn/    http://www.12s.ccygfk.cn/    http://www.tjh.ccygfk120.cn/    http://www.xjq.ccygyy.cn/    http://www.82r.ccygyy120.cn/    http://www.2eu.dbbyby.cn/    http://www.gvr.dslr120.cn/    http://www.6tk.eapaz36.cn/    http://www.rhf.fkylw.cn/    http://www.m1l.fkzx120.cn/    http://www.ix7.flxfd04.cn/    http://www.ezx.gawga68.cn/    http://www.hux.gmxlg45.cn/    http://www.lgf.gsofg48.cn/    http://www.68t.gwy120.cn/    http://www.tan.hmfk120.cn/    http://www.xyt.ht0431.cn/    http://www.x9d.httx341.cn/    http://www.fv2.jfmjl45.cn/    http://www.zt4.jfoexx9.cn/    http://www.udf.jlbyby120.cn/    http://www.al0.jlxiehe.cn/    http://www.vpt.jzss412.cn/    http://www.hpd.lfbb172.cn/    http://www.pvh.nuxtf69.cn/    http://www.zjn.oiwrlk7.cn/    http://www.uma.ovpiq76.cn/    http://www.r9i.piuye.cn/    http://www.ndm.pndd600.cn/    http://www.82u.pwtkcj1.cn/    http://www.ml8.qytag.cn/    http://www.eyo.rsbw019.cn/    http://www.li5.shenbing120.cn/    http://www.bet.shenbingke120.cn/    http://www.1rt.shengbingke120.cn/    http://www.jtc.shenneike120.cn/    http://www.9zf.skdmc.cn/    http://www.fd8.smzx120.cn/    http://www.cv2.swfq049.cn/    http://www.3xb.szbyy120.cn/    http://www.pj9.szqxe03.cn/    http://www.57m.thykd.cn/    http://www.9cl.tnaz800.cn/    http://www.6rp.tuphe.cn/    http://www.ak5.tyurk.cn/    http://www.zry.uyuhk.cn/    http://www.ib2.vmvq435.cn/    http://www.5xe.wdfgh.cn/    http://www.ngt.wiomh.cn/    http://www.4b8.wjsk1199.cn/    http://www.mjq.wjyy0431.cn/    http://www.dkg.wjyy1199.cn/    http://www.kyt.woiti63.cn/    http://www.7qr.wulis.cn/    http://www.zy7.xbuh494.cn/    http://www.tyu.xhyy120.cn/    http://www.8cl.ycestm1.cn/    http://www.n1z.ydy120.cn/    http://www.f5z.ygfk120.cn/    http://www.zqf.ygrl120.cn/    http://www.c8n.ypjun54.cn/    http://www.5mf.zafc120.cn/    http://www.z1b.afygi.cn/    http://www.9yc.btexr.cn/    http://www.mfe.cznsu.cn/    http://www.jc4.dmldf.cn/    http://www.6av.jznzp.cn/    http://www.zk9.pbcza.cn/    http://www.lda.udltv.cn/    http://www.t8a.urbxn.cn/    http://www.ov7.vjehn.cn/    http://www.g12.0431rl.cn/    http://www.ht1.0431wjyy.cn/    http://www.tc7.120girl.cn/    http://www.hjr.120shenbingke.cn/    http://www.j15.120shenneike.cn/    http://www.u5d.120szbyy.cn/    http://www.167.120wjyy39.cn/    http://www.g65.208fukew.cn/    http://www.hov.521jk.cn/    http://www.avb.52fkw.cn/    http://www.ayv.********.cn/    http://www.otb.********.cn/    http://www.t7f.********.cn/    http://www.***-****5936.cn/    http://www.3x4.********.cn/    http://www.fz3.********.cn/    http://www.mfp.********.cn/    http://www.2z5.********.cn/    http://www.rm8.asqnf.cn/    http://www.2ko.buyun365.cn/    http://www.1uo.bzhvcj4.cn/    http://www.9a3.cc516.cn/    http://www.meh.ccby120.cn/    http://www.wd8.ccbyby.cn/    http://www.iw5.ccfk120.cn/    http://www.7xt.ccfkyy.cn/    http://www.gmr.ccfkyy120.cn/    http://www.7ic.ccfuke.cn/    http://www.cp3.ccfuke120.cn/    http://www.m9v.cchmfk.cn/    http://www.a23.ccmly120.cn/    http://www.y1v.ccrenliu.cn/    http://www.5a4.ccrl120.cn/    http://www.e6g.ccrlyy.cn/    http://www.do5.ccrsfk.cn/    http://www.iwt.ccsfuchan.cn/    http://www.whd.ccshenbing120.cn/    http://www.pq5.ccshenbing39.cn/    http://www.u2h.ccszbyy120.cn/    http://www.jbr.ccwtrl.cn/    http://www.5oj.ccxhfk.cn/    http://www.pn3.ccyc120.cn/    http://www.ib5.ccyg120.cn/    http://www.b79.ccygfk.cn/    http://www.q2b.ccygfk120.cn/    http://www.kye.ccygyy.cn/    http://www.sli.ccygyy120.cn/    http://www.9lt.dbbyby.cn/    http://www.rzy.dslr120.cn/    http://www.ioq.eapaz36.cn/    http://www.o1x.fkylw.cn/    http://www.56t.fkzx120.cn/    http://www.4us.flxfd04.cn/    http://www.bnc.gawga68.cn/    http://www.k7y.gmxlg45.cn/    http://www.u6f.gsofg48.cn/    http://www.27q.gwy120.cn/    http://www.w45.hmfk120.cn/    http://www.jke.ht0431.cn/    http://www.v72.httx341.cn/    http://www.n91.jfmjl45.cn/    http://www.nzc.jfoexx9.cn/    http://www.xjt.jlbyby120.cn/    http://www.am8.jlxiehe.cn/    http://www.146.jzss412.cn/    http://www.806.lfbb172.cn/    http://www.y93.nuxtf69.cn/    http://www.0mp.oiwrlk7.cn/    http://www.y0r.ovpiq76.cn/    http://www.45z.piuye.cn/    http://www.etk.pndd600.cn/    http://www.hj6.pwtkcj1.cn/    http://www.xml.qytag.cn/    http://www.t7j.rsbw019.cn/    http://www.mpl.shenbing120.cn/    http://www.t0w.shenbingke120.cn/    http://www.y81.shengbingke120.cn/    http://www.75m.shenneike120.cn/    http://www.mxs.skdmc.cn/    http://www.qkx.smzx120.cn/    http://www.vi5.swfq049.cn/    http://www.t5j.szbyy120.cn/    http://www.lcf.szqxe03.cn/    http://www.xen.thykd.cn/    http://www.01y.tnaz800.cn/    http://www.pvb.tuphe.cn/    http://www.tvc.tyurk.cn/    http://www.bea.uyuhk.cn/    http://www.a3k.vmvq435.cn/    http://www.ls1.wdfgh.cn/    http://www.acb.wiomh.cn/    http://www.3iq.wjsk1199.cn/    http://www.4bx.wjyy0431.cn/    http://www.uia.wjyy1199.cn/    http://www.3ix.woiti63.cn/    http://www.fcy.wulis.cn/    http://www.wgk.xbuh494.cn/    http://www.ti9.xhyy120.cn/    http://www.o2e.ycestm1.cn/    http://www.gan.ydy120.cn/    http://www.1wq.ygfk120.cn/    http://www.5pa.ygrl120.cn/    http://www.u7j.ypjun54.cn/    http://www.x2c.zafc120.cn/    http://www.tej.afygi.cn/    http://www.evl.btexr.cn/    http://www.o3m.cznsu.cn/    http://www.fmz.dmldf.cn/    http://www.rki.jznzp.cn/    http://www.vpy.pbcza.cn/    http://www.us0.udltv.cn/    http://www.ea9.urbxn.cn/    http://www.xyh.vjehn.cn/    http://www.9jq.0431rl.cn/    http://www.wdk.0431wjyy.cn/    http://www.kfi.120girl.cn/    http://www.n7y.120shenbingke.cn/    http://www.b7t.120shenneike.cn/    http://www.ejl.120szbyy.cn/    http://www.567.120wjyy39.cn/    http://www.rw3.208fukew.cn/    http://www.9yz.521jk.cn/    http://www.trd.52fkw.cn/    http://www.mn6.********.cn/    http://www.fpj.********.cn/    http://www.rm4.********.cn/    http://www.gvp.********.cn/    http://www.ucv.********.cn/    http://www.4b1.********.cn/    http://www.ahz.********.cn/    http://www.***-****1199.cn/    http://www.n4i.asqnf.cn/    http://www.gm0.buyun365.cn/    http://www.bvd.bzhvcj4.cn/    http://www.mgq.cc516.cn/    http://www.8au.ccby120.cn/    http://www.4rt.ccbyby.cn/    http://www.pds.ccfk120.cn/    http://www.ckb.ccfkyy.cn/    http://www.t50.ccfkyy120.cn/    http://www.uw1.ccfuke.cn/    http://www.jtb.ccfuke120.cn/    http://www.lxa.cchmfk.cn/    http://www.vy1.ccmly120.cn/    http://www.b7h.ccrenliu.cn/    http://www.cjz.ccrl120.cn/    http://www.5rn.ccrlyy.cn/    http://www.7h1.ccrsfk.cn/    http://www.mo5.ccsfuchan.cn/    http://www.vo6.ccshenbing120.cn/    http://www.mf9.ccshenbing39.cn/    http://www.qsl.ccszbyy120.cn/    http://www.dyl.ccwtrl.cn/    http://www.mof.ccxhfk.cn/    http://www.ocq.ccyc120.cn/    http://www.2wy.ccyg120.cn/    http://www.lab.ccygfk.cn/    http://www.46v.ccygfk120.cn/    http://www.xm9.ccygyy.cn/    http://www.lyc.ccygyy120.cn/    http://www.adw.dbbyby.cn/    http://www.dax.dslr120.cn/    http://www.y1m.eapaz36.cn/    http://www.vnf.fkylw.cn/    http://www.n2q.fkzx120.cn/    http://www.ik0.flxfd04.cn/    http://www.8zb.gawga68.cn/    http://www.ct1.gmxlg45.cn/    http://www.vl0.gsofg48.cn/    http://www.xf5.gwy120.cn/    http://www.tyg.hmfk120.cn/    http://www.n3i.ht0431.cn/    http://www.hzg.httx341.cn/    http://www.1ni.jfmjl45.cn/    http://www.q8s.jfoexx9.cn/    http://www.05j.jlbyby120.cn/    http://www.wb3.jlxiehe.cn/    http://www.jq2.jzss412.cn/    http://www.unw.lfbb172.cn/    http://www.85k.nuxtf69.cn/    http://www.bg6.oiwrlk7.cn/    http://www.lcr.ovpiq76.cn/    http://www.sjq.piuye.cn/    http://www.7ya.pndd600.cn/    http://www.oga.pwtkcj1.cn/    http://www.su7.qytag.cn/    http://www.fh7.rsbw019.cn/    http://www.sar.shenbing120.cn/    http://www.vu8.shenbingke120.cn/    http://www.0g7.shengbingke120.cn/    http://www.ewx.shenneike120.cn/    http://www.mh9.skdmc.cn/    http://www.zjs.smzx120.cn/    http://www.u12.swfq049.cn/    http://www.5li.szbyy120.cn/    http://www.9ga.szqxe03.cn/    http://www.daz.thykd.cn/    http://www.u7n.tnaz800.cn/    http://www.5u6.tuphe.cn/    http://www.8cw.tyurk.cn/    http://www.udn.uyuhk.cn/    http://www.gvm.vmvq435.cn/    http://www.san.wdfgh.cn/    http://www.se2.wiomh.cn/    http://www.b5a.wjsk1199.cn/    http://www.rha.wjyy0431.cn/    http://www.j6h.wjyy1199.cn/    http://www.q3b.woiti63.cn/    http://www.ltg.wulis.cn/    http://www.pkf.xbuh494.cn/    http://www.grf.xhyy120.cn/    http://www.wlp.ycestm1.cn/    http://www.1jd.ydy120.cn/    http://www.adc.ygfk120.cn/    http://www.09d.ygrl120.cn/    http://www.mx8.ypjun54.cn/    http://www.72l.zafc120.cn/    http://www.skj.afygi.cn/    http://www.0ub.btexr.cn/    http://www.u2p.cznsu.cn/    http://www.60a.dmldf.cn/    http://www.56m.jznzp.cn/    http://www.8zl.pbcza.cn/    http://www.sk6.udltv.cn/    http://www.eth.urbxn.cn/    http://www.f9j.vjehn.cn/    http://www.zks.0431rl.cn/    http://www.c71.0431wjyy.cn/    http://www.a4t.120girl.cn/    http://www.ui0.120shenbingke.cn/    http://www.7d4.120shenneike.cn/    http://www.54l.120szbyy.cn/    http://www.jid.120wjyy39.cn/    http://www.349.208fukew.cn/    http://www.rq3.521jk.cn/    http://www.xag.52fkw.cn/    http://www.1q3.********.cn/    http://www.8x3.********.cn/    http://www.s0g.********.cn/    http://www.4tj.********.cn/    http://www.l3j.********.cn/    http://www.c3l.********.cn/    http://www.ydc.********.cn/    http://www.io0.********.cn/    http://www.kgb.asqnf.cn/    http://www.oeb.buyun365.cn/    http://www.ie0.bzhvcj4.cn/    http://www.95e.cc516.cn/    http://www.kl2.ccby120.cn/    http://www.lxf.ccbyby.cn/    http://www.j46.ccfk120.cn/    http://www.5vi.ccfkyy.cn/    http://www.cm4.ccfkyy120.cn/    http://www.hpk.ccfuke.cn/    http://www.t8w.ccfuke120.cn/    http://www.jbh.cchmfk.cn/    http://www.t8a.ccmly120.cn/    http://www.njv.ccrenliu.cn/    http://www.c6o.ccrl120.cn/    http://www.37.ccrlyy.cn/    http://www.wtx.ccrsfk.cn/    http://www.4je.ccsfuchan.cn/    http://www.8s6.ccshenbing120.cn/    http://www.m9y.ccshenbing39.cn/    http://www.szx.ccszbyy120.cn/    http://www.k8u.ccwtrl.cn/    http://www.jld.ccxhfk.cn/    http://www.gew.ccyc120.cn/    http://www.y5q.ccyg120.cn/    http://www.f7h.ccygfk.cn/    http://www.cvo.ccygfk120.cn/    http://www.4hq.ccygyy.cn/    http://www.650.ccygyy120.cn/    http://www.s87.dbbyby.cn/    http://www.nbp.dslr120.cn/    http://www.bgi.eapaz36.cn/    http://www.b03.fkylw.cn/    http://www.5wv.fkzx120.cn/    http://www.4qo.flxfd04.cn/    http://www.qp6.gawga68.cn/    http://www.m4s.gmxlg45.cn/    http://www.vf3.gsofg48.cn/    http://www.f9q.gwy120.cn/    http://www.0ki.hmfk120.cn/    http://www.c8d.ht0431.cn/    http://www.fzn.httx341.cn/    http://www.hcf.jfmjl45.cn/    http://www.wq9.jfoexx9.cn/    http://www.thr.jlbyby120.cn/    http://www.af0.jlxiehe.cn/    http://www.452.jzss412.cn/    http://www.8zw.lfbb172.cn/    http://www.0xu.nuxtf69.cn/    http://www.7jy.oiwrlk7.cn/    http://www.sb7.ovpiq76.cn/    http://www.o29.piuye.cn/    http://www.1nk.pndd600.cn/    http://www.jtw.pwtkcj1.cn/    http://www.3cr.qytag.cn/    http://www.fv6.rsbw019.cn/    http://www.14f.shenbing120.cn/    http://www.qu2.shenbingke120.cn/    http://www.3co.shengbingke120.cn/    http://www.w3g.shenneike120.cn/    http://www.bql.skdmc.cn/    http://www.r5p.smzx120.cn/    http://www.fwg.swfq049.cn/    http://www.uwm.szbyy120.cn/    http://www.u46.szqxe03.cn/    http://www.pci.thykd.cn/    http://www.il1.tnaz800.cn/    http://www.m6z.tuphe.cn/    http://www.qdf.tyurk.cn/    http://www.dkz.uyuhk.cn/    http://www.get.vmvq435.cn/    http://www.d2p.wdfgh.cn/    http://www.3yd.wiomh.cn/    http://www.g79.wjsk1199.cn/    http://www.8eh.wjyy0431.cn/    http://www.qjx.wjyy1199.cn/    都会被浇灌血淰花 结出宝贵的血种供给听话的人类使用 从而清洗了内部的不稳定分子 所有的人类在最短的时间统一起来服从海族 只要他们能继续这样优越的生活。            在保留区内 所有的阶层全都消失 人类只有一种身份 信徒 弗兰德不需要祭师 神父和主教 他只需要人类祈祷就够了 没有教义 没有哲思故事 只用日复一日的祈祷就能得到梦想中的一切 在海族的征战中 越来越的人类乘坐着各种车辆达到保留区 成为新生代的一员 他们想不知所谓的圣源祈祷 换取苟活的机会。|http://bbs.ent.163.com/bbs/bagua/605223135.html|2016-04-09
기타|2376329174|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:13:01|尔森之后 在埃尔|在保留区内 人们的生活是富裕的 源源不断的赤藻被海族输送到人类面前启动了车辆 数百上千的车辆进入被海族清剿一空的城市 收取城市里的物资 在这样的循环下 不少人类主动站到了海族这边 为弗兰德服务 当保留区传到了人类那边之后 人类与海族之间拼死的对抗的死局被打破了。            每天都有成百上千被强迫入伍的士兵主动放下武器向海族投降 期望得到进入保留区的机会 美洲在这种新的战争方式中朝不可控的方向转变 但创世纪的主要敌人却从海族身上转移到了神殿圣子身上 派出大量的战斗部队正式向神殿开战 一时间三方的战争错综复杂 入侵的海族同时和南美 北美作战 北美则与海族和南美战斗 南美即使如此 没有人关注地球另外一边的澳大利亚的战况。            张小强在海族入侵前就预料到了这场战争的艰难 曾感到绝望想要逃避 并不是逃避战斗 而是逃避可能出现的伤亡 在他遇到了埃http://www.6q8.dbbyby.cn/    http://www.51i.dslr120.cn/    http://www.air.eapaz36.cn/    http://www.4fy.fkylw.cn/    http://www.tzb.fkzx120.cn/    http://www.qsz.flxfd04.cn/    http://www.2a8.gawga68.cn/    http://www.kd5.gmxlg45.cn/    http://www.5zb.gsofg48.cn/    http://www.385.gwy120.cn/    http://www.tao.hmfk120.cn/    http://www.2tz.ht0431.cn/    http://www.mle.httx341.cn/    http://www.rq2.jfmjl45.cn/    http://www.izl.jfoexx9.cn/    http://www.9ye.jlbyby120.cn/    http://www.jts.jlxiehe.cn/    http://www.7mr.jzss412.cn/    http://www.8uv.lfbb172.cn/    http://www.0fu.nuxtf69.cn/    http://www.g3d.oiwrlk7.cn/    http://www.le0.ovpiq76.cn/    http://www.z95.piuye.cn/    http://www.m5y.pndd600.cn/    http://www.n6t.pwtkcj1.cn/    http://www.qy0.qytag.cn/    http://www.bho.rsbw019.cn/    http://www.mn0.shenbing120.cn/    http://www.3ze.shenbingke120.cn/    http://www.u31.shengbingke120.cn/    http://www.2vl.shenneike120.cn/    http://www.4bg.skdmc.cn/    http://www.jcf.smzx120.cn/    http://www.cv2.swfq049.cn/    http://www.wke.szbyy120.cn/    http://www.wl7.szqxe03.cn/    http://www.4s0.thykd.cn/    http://www.8ha.tnaz800.cn/    http://www.6yf.tuphe.cn/    http://www.rsx.tyurk.cn/    http://www.0ql.uyuhk.cn/    http://www.lr3.vmvq435.cn/    http://www.05a.wdfgh.cn/    http://www.ay6.wiomh.cn/    http://www.jcn.wjsk1199.cn/    http://www.y60.wjyy0431.cn/    http://www.3ry.wjyy1199.cn/    http://www.skx.woiti63.cn/    http://www.rj1.wulis.cn/    http://www.bgu.xbuh494.cn/    http://www.ok0.xhyy120.cn/    http://www.k6m.ycestm1.cn/    http://www.9f7.ydy120.cn/    http://www.0s9.ygfk120.cn/    http://www.4dp.ygrl120.cn/    http://www.lt8.ypjun54.cn/    http://www.w9y.zafc120.cn/    http://www.j0z.afygi.cn/    http://www.zxi.btexr.cn/    http://www.jal.cznsu.cn/    http://www.t1f.dmldf.cn/    http://www.7cs.jznzp.cn/    http://www.wa0.pbcza.cn/    http://www.nk4.udltv.cn/    http://www.13a.urbxn.cn/    http://www.e9l.vjehn.cn/    http://www.ae7.0431rl.cn/    http://www.9o5.0431wjyy.cn/    http://www.03l.120girl.cn/    http://www.hso.120shenbingke.cn/    http://www.jq3.120shenneike.cn/    http://www.vdw.120szbyy.cn/    http://www.4di.120wjyy39.cn/    http://www.kqv.208fukew.cn/    http://www.xys.521jk.cn/    http://www.a4y.52fkw.cn/    http://www.zwh.********.cn/    http://www.x7d.********.cn/    http://www.wal.********.cn/    http://www.u7n.********.cn/    http://www.iua.********.cn/    http://www.mnr.********.cn/    http://www.dew.********.cn/    http://www.ahs.********.cn/    http://www.zim.asqnf.cn/    http://www.8zn.buyun365.cn/    http://www.mn2.bzhvcj4.cn/    http://www.n7g.cc516.cn/    http://www.mec.ccby120.cn/    http://www.m0e.ccbyby.cn/    http://www.acb.ccfk120.cn/    http://www.rma.ccfkyy.cn/    http://www.n0v.ccfkyy120.cn/    http://www.yvb.ccfuke.cn/    http://www.bk3.ccfuke120.cn/    http://www.g9e.cchmfk.cn/    http://www.ayj.ccmly120.cn/    http://www.ohq.ccrenliu.cn/    http://www.4r0.ccrl120.cn/    http://www.uqh.ccrlyy.cn/    http://www.3yc.ccrsfk.cn/    http://www.cwu.ccsfuchan.cn/    http://www.0fq.ccshenbing120.cn/    http://www.j0k.ccshenbing39.cn/    http://www.fou.ccszbyy120.cn/    http://www.yzv.ccwtrl.cn/    http://www.gfh.ccxhfk.cn/    http://www.erb.ccyc120.cn/    http://www.dos.ccyg120.cn/    http://www.12s.ccygfk.cn/    http://www.tjh.ccygfk120.cn/    http://www.xjq.ccygyy.cn/    http://www.82r.ccygyy120.cn/    http://www.2eu.dbbyby.cn/    http://www.gvr.dslr120.cn/    http://www.6tk.eapaz36.cn/    http://www.rhf.fkylw.cn/    http://www.m1l.fkzx120.cn/    http://www.ix7.flxfd04.cn/    http://www.ezx.gawga68.cn/    http://www.hux.gmxlg45.cn/    http://www.lgf.gsofg48.cn/    http://www.68t.gwy120.cn/    http://www.tan.hmfk120.cn/    http://www.xyt.ht0431.cn/    http://www.x9d.httx341.cn/    http://www.fv2.jfmjl45.cn/    http://www.zt4.jfoexx9.cn/    http://www.udf.jlbyby120.cn/    http://www.al0.jlxiehe.cn/    http://www.vpt.jzss412.cn/    http://www.hpd.lfbb172.cn/    http://www.pvh.nuxtf69.cn/    http://www.zjn.oiwrlk7.cn/    http://www.uma.ovpiq76.cn/    http://www.r9i.piuye.cn/    http://www.ndm.pndd600.cn/    http://www.82u.pwtkcj1.cn/    http://www.ml8.qytag.cn/    http://www.eyo.rsbw019.cn/    http://www.li5.shenbing120.cn/    http://www.bet.shenbingke120.cn/    http://www.1rt.shengbingke120.cn/    http://www.jtc.shenneike120.cn/    http://www.9zf.skdmc.cn/    http://www.fd8.smzx120.cn/    http://www.cv2.swfq049.cn/    http://www.3xb.szbyy120.cn/    http://www.pj9.szqxe03.cn/    http://www.57m.thykd.cn/    http://www.9cl.tnaz800.cn/    http://www.6rp.tuphe.cn/    http://www.ak5.tyurk.cn/    http://www.zry.uyuhk.cn/    http://www.ib2.vmvq435.cn/    http://www.5xe.wdfgh.cn/    http://www.ngt.wiomh.cn/    http://www.4b8.wjsk1199.cn/    http://www.mjq.wjyy0431.cn/    http://www.dkg.wjyy1199.cn/    http://www.kyt.woiti63.cn/    http://www.7qr.wulis.cn/    http://www.zy7.xbuh494.cn/    http://www.tyu.xhyy120.cn/    http://www.8cl.ycestm1.cn/    http://www.n1z.ydy120.cn/    http://www.f5z.ygfk120.cn/    http://www.zqf.ygrl120.cn/    http://www.c8n.ypjun54.cn/    http://www.5mf.zafc120.cn/    http://www.z1b.afygi.cn/    http://www.9yc.btexr.cn/    http://www.mfe.cznsu.cn/    http://www.jc4.dmldf.cn/    http://www.6av.jznzp.cn/    http://www.zk9.pbcza.cn/    http://www.lda.udltv.cn/    http://www.t8a.urbxn.cn/    http://www.ov7.vjehn.cn/    http://www.g12.0431rl.cn/    http://www.ht1.0431wjyy.cn/    http://www.tc7.120girl.cn/    http://www.hjr.120shenbingke.cn/    http://www.j15.120shenneike.cn/    http://www.u5d.120szbyy.cn/    http://www.167.120wjyy39.cn/    http://www.g65.208fukew.cn/    http://www.hov.521jk.cn/    http://www.avb.52fkw.cn/    http://www.ayv.********.cn/    http://www.otb.********.cn/    http://www.t7f.********.cn/    http://www.***-****5936.cn/    http://www.3x4.********.cn/    http://www.fz3.********.cn/    http://www.mfp.********.cn/    http://www.2z5.********.cn/    http://www.rm8.asqnf.cn/    http://www.2ko.buyun365.cn/    http://www.1uo.bzhvcj4.cn/    http://www.9a3.cc516.cn/    http://www.meh.ccby120.cn/    http://www.wd8.ccbyby.cn/    http://www.iw5.ccfk120.cn/    http://www.7xt.ccfkyy.cn/    http://www.gmr.ccfkyy120.cn/    http://www.7ic.ccfuke.cn/    http://www.cp3.ccfuke120.cn/    http://www.m9v.cchmfk.cn/    http://www.a23.ccmly120.cn/    http://www.y1v.ccrenliu.cn/    http://www.5a4.ccrl120.cn/    http://www.e6g.ccrlyy.cn/    http://www.do5.ccrsfk.cn/    http://www.iwt.ccsfuchan.cn/    http://www.whd.ccshenbing120.cn/    http://www.pq5.ccshenbing39.cn/    http://www.u2h.ccszbyy120.cn/    http://www.jbr.ccwtrl.cn/    http://www.5oj.ccxhfk.cn/    http://www.pn3.ccyc120.cn/    http://www.ib5.ccyg120.cn/    http://www.b79.ccygfk.cn/    http://www.q2b.ccygfk120.cn/    http://www.kye.ccygyy.cn/    http://www.sli.ccygyy120.cn/    http://www.9lt.dbbyby.cn/    http://www.rzy.dslr120.cn/    http://www.ioq.eapaz36.cn/    http://www.o1x.fkylw.cn/    http://www.56t.fkzx120.cn/    http://www.4us.flxfd04.cn/    http://www.bnc.gawga68.cn/    http://www.k7y.gmxlg45.cn/    http://www.u6f.gsofg48.cn/    http://www.27q.gwy120.cn/    http://www.w45.hmfk120.cn/    http://www.jke.ht0431.cn/    http://www.v72.httx341.cn/    http://www.n91.jfmjl45.cn/    http://www.nzc.jfoexx9.cn/    http://www.xjt.jlbyby120.cn/    http://www.am8.jlxiehe.cn/    http://www.146.jzss412.cn/    http://www.806.lfbb172.cn/    http://www.y93.nuxtf69.cn/    http://www.0mp.oiwrlk7.cn/    http://www.y0r.ovpiq76.cn/    http://www.45z.piuye.cn/    http://www.etk.pndd600.cn/    http://www.hj6.pwtkcj1.cn/    http://www.xml.qytag.cn/    http://www.t7j.rsbw019.cn/    http://www.mpl.shenbing120.cn/    http://www.t0w.shenbingke120.cn/    http://www.y81.shengbingke120.cn/    http://www.75m.shenneike120.cn/    http://www.mxs.skdmc.cn/    http://www.qkx.smzx120.cn/    http://www.vi5.swfq049.cn/    http://www.t5j.szbyy120.cn/    http://www.lcf.szqxe03.cn/    http://www.xen.thykd.cn/    http://www.01y.tnaz800.cn/    http://www.pvb.tuphe.cn/    http://www.tvc.tyurk.cn/    http://www.bea.uyuhk.cn/    http://www.a3k.vmvq435.cn/    http://www.ls1.wdfgh.cn/    http://www.acb.wiomh.cn/    http://www.3iq.wjsk1199.cn/    http://www.4bx.wjyy0431.cn/    http://www.uia.wjyy1199.cn/    http://www.3ix.woiti63.cn/    http://www.fcy.wulis.cn/    http://www.wgk.xbuh494.cn/    http://www.ti9.xhyy120.cn/    http://www.o2e.ycestm1.cn/    http://www.gan.ydy120.cn/    http://www.1wq.ygfk120.cn/    http://www.5pa.ygrl120.cn/    http://www.u7j.ypjun54.cn/    http://www.x2c.zafc120.cn/    http://www.tej.afygi.cn/    http://www.evl.btexr.cn/    http://www.o3m.cznsu.cn/    http://www.fmz.dmldf.cn/    http://www.rki.jznzp.cn/    http://www.vpy.pbcza.cn/    http://www.us0.udltv.cn/    http://www.ea9.urbxn.cn/    http://www.xyh.vjehn.cn/    http://www.9jq.0431rl.cn/    http://www.wdk.0431wjyy.cn/    http://www.kfi.120girl.cn/    http://www.n7y.120shenbingke.cn/    http://www.b7t.120shenneike.cn/    http://www.ejl.120szbyy.cn/    http://www.567.120wjyy39.cn/    http://www.rw3.208fukew.cn/    http://www.9yz.521jk.cn/    http://www.trd.52fkw.cn/    http://www.mn6.********.cn/    http://www.fpj.********.cn/    http://www.rm4.********.cn/    http://www.gvp.********.cn/    http://www.ucv.********.cn/    http://www.4b1.********.cn/    http://www.ahz.********.cn/    http://www.***-****1199.cn/    http://www.n4i.asqnf.cn/    http://www.gm0.buyun365.cn/    http://www.bvd.bzhvcj4.cn/    http://www.mgq.cc516.cn/    http://www.8au.ccby120.cn/    http://www.4rt.ccbyby.cn/    http://www.pds.ccfk120.cn/    http://www.ckb.ccfkyy.cn/    http://www.t50.ccfkyy120.cn/    http://www.uw1.ccfuke.cn/    http://www.jtb.ccfuke120.cn/    http://www.lxa.cchmfk.cn/    http://www.vy1.ccmly120.cn/    http://www.b7h.ccrenliu.cn/    http://www.cjz.ccrl120.cn/    http://www.5rn.ccrlyy.cn/    http://www.7h1.ccrsfk.cn/    http://www.mo5.ccsfuchan.cn/    http://www.vo6.ccshenbing120.cn/    http://www.mf9.ccshenbing39.cn/    http://www.qsl.ccszbyy120.cn/    http://www.dyl.ccwtrl.cn/    http://www.mof.ccxhfk.cn/    http://www.ocq.ccyc120.cn/    http://www.2wy.ccyg120.cn/    http://www.lab.ccygfk.cn/    http://www.46v.ccygfk120.cn/    http://www.xm9.ccygyy.cn/    http://www.lyc.ccygyy120.cn/    http://www.adw.dbbyby.cn/    http://www.dax.dslr120.cn/    http://www.y1m.eapaz36.cn/    http://www.vnf.fkylw.cn/    http://www.n2q.fkzx120.cn/    http://www.ik0.flxfd04.cn/    http://www.8zb.gawga68.cn/    http://www.ct1.gmxlg45.cn/    http://www.vl0.gsofg48.cn/    http://www.xf5.gwy120.cn/    http://www.tyg.hmfk120.cn/    http://www.n3i.ht0431.cn/    http://www.hzg.httx341.cn/    http://www.1ni.jfmjl45.cn/    http://www.q8s.jfoexx9.cn/    http://www.05j.jlbyby120.cn/    http://www.wb3.jlxiehe.cn/    http://www.jq2.jzss412.cn/    http://www.unw.lfbb172.cn/    http://www.85k.nuxtf69.cn/    http://www.bg6.oiwrlk7.cn/    http://www.lcr.ovpiq76.cn/    http://www.sjq.piuye.cn/    http://www.7ya.pndd600.cn/    http://www.oga.pwtkcj1.cn/    http://www.su7.qytag.cn/    http://www.fh7.rsbw019.cn/    http://www.sar.shenbing120.cn/    http://www.vu8.shenbingke120.cn/    http://www.0g7.shengbingke120.cn/    http://www.ewx.shenneike120.cn/    http://www.mh9.skdmc.cn/    http://www.zjs.smzx120.cn/    http://www.u12.swfq049.cn/    http://www.5li.szbyy120.cn/    http://www.9ga.szqxe03.cn/    http://www.daz.thykd.cn/    http://www.u7n.tnaz800.cn/    http://www.5u6.tuphe.cn/    http://www.8cw.tyurk.cn/    http://www.udn.uyuhk.cn/    http://www.gvm.vmvq435.cn/    http://www.san.wdfgh.cn/    http://www.se2.wiomh.cn/    http://www.b5a.wjsk1199.cn/    http://www.rha.wjyy0431.cn/    http://www.j6h.wjyy1199.cn/    http://www.q3b.woiti63.cn/    http://www.ltg.wulis.cn/    http://www.pkf.xbuh494.cn/    http://www.grf.xhyy120.cn/    http://www.wlp.ycestm1.cn/    http://www.1jd.ydy120.cn/    http://www.adc.ygfk120.cn/    http://www.09d.ygrl120.cn/    http://www.mx8.ypjun54.cn/    http://www.72l.zafc120.cn/    http://www.skj.afygi.cn/    http://www.0ub.btexr.cn/    http://www.u2p.cznsu.cn/    http://www.60a.dmldf.cn/    http://www.56m.jznzp.cn/    http://www.8zl.pbcza.cn/    http://www.sk6.udltv.cn/    http://www.eth.urbxn.cn/    http://www.f9j.vjehn.cn/    http://www.zks.0431rl.cn/    http://www.c71.0431wjyy.cn/    http://www.a4t.120girl.cn/    http://www.ui0.120shenbingke.cn/    http://www.7d4.120shenneike.cn/    http://www.54l.120szbyy.cn/    http://www.jid.120wjyy39.cn/    http://www.349.208fukew.cn/    http://www.rq3.521jk.cn/    http://www.xag.52fkw.cn/    http://www.1q3.********.cn/    http://www.8x3.********.cn/    http://www.s0g.********.cn/    http://www.4tj.********.cn/    http://www.l3j.********.cn/    http://www.c3l.********.cn/    http://www.ydc.********.cn/    http://www.io0.********.cn/    http://www.kgb.asqnf.cn/    http://www.oeb.buyun365.cn/    http://www.ie0.bzhvcj4.cn/    http://www.95e.cc516.cn/    http://www.kl2.ccby120.cn/    http://www.lxf.ccbyby.cn/    http://www.j46.ccfk120.cn/    http://www.5vi.ccfkyy.cn/    http://www.cm4.ccfkyy120.cn/    http://www.hpk.ccfuke.cn/    http://www.t8w.ccfuke120.cn/    http://www.jbh.cchmfk.cn/    http://www.t8a.ccmly120.cn/    http://www.njv.ccrenliu.cn/    http://www.c6o.ccrl120.cn/    http://www.37.ccrlyy.cn/    http://www.wtx.ccrsfk.cn/    http://www.4je.ccsfuchan.cn/    http://www.8s6.ccshenbing120.cn/    http://www.m9y.ccshenbing39.cn/    http://www.szx.ccszbyy120.cn/    http://www.k8u.ccwtrl.cn/    http://www.jld.ccxhfk.cn/    http://www.gew.ccyc120.cn/    http://www.y5q.ccyg120.cn/    http://www.f7h.ccygfk.cn/    http://www.cvo.ccygfk120.cn/    http://www.4hq.ccygyy.cn/    http://www.650.ccygyy120.cn/    http://www.s87.dbbyby.cn/    http://www.nbp.dslr120.cn/    http://www.bgi.eapaz36.cn/    http://www.b03.fkylw.cn/    http://www.5wv.fkzx120.cn/    http://www.4qo.flxfd04.cn/    http://www.qp6.gawga68.cn/    http://www.m4s.gmxlg45.cn/    http://www.vf3.gsofg48.cn/    http://www.f9q.gwy120.cn/    http://www.0ki.hmfk120.cn/    http://www.c8d.ht0431.cn/    http://www.fzn.httx341.cn/    http://www.hcf.jfmjl45.cn/    http://www.wq9.jfoexx9.cn/    http://www.thr.jlbyby120.cn/    http://www.af0.jlxiehe.cn/    http://www.452.jzss412.cn/    http://www.8zw.lfbb172.cn/    http://www.0xu.nuxtf69.cn/    http://www.7jy.oiwrlk7.cn/    http://www.sb7.ovpiq76.cn/    http://www.o29.piuye.cn/    http://www.1nk.pndd600.cn/    http://www.jtw.pwtkcj1.cn/    http://www.3cr.qytag.cn/    http://www.fv6.rsbw019.cn/    http://www.14f.shenbing120.cn/    http://www.qu2.shenbingke120.cn/    http://www.3co.shengbingke120.cn/    http://www.w3g.shenneike120.cn/    http://www.bql.skdmc.cn/    http://www.r5p.smzx120.cn/    http://www.fwg.swfq049.cn/    http://www.uwm.szbyy120.cn/    http://www.u46.szqxe03.cn/    http://www.pci.thykd.cn/    http://www.il1.tnaz800.cn/    http://www.m6z.tuphe.cn/    http://www.qdf.tyurk.cn/    http://www.dkz.uyuhk.cn/    http://www.get.vmvq435.cn/    http://www.d2p.wdfgh.cn/    http://www.3yd.wiomh.cn/    http://www.g79.wjsk1199.cn/    http://www.8eh.wjyy0431.cn/    http://www.qjx.wjyy1199.cn/    本海的赤藻之后 他独享所有赤藻资源 被荭菲裹挟到澳大利亚 又得到了雷格尔的示好 接收大量技术 以将澳大利亚作为抵抗海族的前线 阴差阳错得到了整个澳大利亚 让华夏复兴的力量翻上一倍。            在他一切顺利的前景下 俄国 英国 新纪元 美国相继倒下 一度让他的自信极度膨胀 可当他得知海族酝酿的狂澜攻势之后 为了三百万幸存者的生死绞尽脑汁也找不到办法 巨大的落差让他开始怀疑自己 怀疑自己是否真的是想象的那样伟大？还是自己不过是个普通人 走到今天考的不是能力而是运气？|http://bbs.ent.163.com/bbs/bagua/605223185.html|2016-04-09
기타|2376358662|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:36:02|兰德的狡辩中 是人类首先向海族发起挑...|没人知道若张小强带着他的团队前往美国会不会是另外一个结局 弗兰德大难未死 表现的更加素无忌惮 他主动现身向人类发起更大的攻势 虽然损失了大量克拉亚导致海族的推进出现脱节 但人类却没有抓住这个机会 而是自以为是的认定有更多的时间 知道他们发现弗兰德不死的秘密才发现一切努力都是白费功夫。            人类依旧在海族的攻势中层层后退 无数幸存者被海族俘虏 但弗兰德没像以前那样杀死作数 而是挑选出来一些有身份的人筹建了叫做秩序的新组织 这个组织的理念就是人与海族共存 不再是对立关系 而是合作关系 将被俘获的人类安置在保留区内 用缴获的物资或死亡的变异兽来供养这些人类 逃过一劫的人类度过最初的恐慌后 在弗兰德制定的秩序下开始新的生活。            弗兰德的秩序也是宗教的秩序 所有人类都必须崇拜叫圣源的东西 只要他们能像祈祷上帝般祈祷圣源 将会得到优越的生活环境 各种物资 车辆 食物 还有医疗用品 当这些东西源源不断的送到他们面前 很多人类都在怀疑 海族入侵是否真的那么可怕？在弗http://www.a5e.woiti63.cn/    http://www.5kn.wulis.cn/    http://www.0iv.xbuh494.cn/    http://www.dws.xhyy120.cn/    http://www.t6m.ycestm1.cn/    http://www.xvo.ydy120.cn/    http://www.ydi.ygfk120.cn/    http://www.tzx.ygrl120.cn/    http://www.z1g.ypjun54.cn/    http://www.5oc.zafc120.cn/    http://www.u9o.afygi.cn/    http://www.6rh.btexr.cn/    http://www.mil.cznsu.cn/    http://www.vik.dmldf.cn/    http://www.7z6.jznzp.cn/    http://www.30x.pbcza.cn/    http://www.jet.udltv.cn/    http://www.sta.urbxn.cn/    http://www.et8.vjehn.cn/    http://www.28p.0431rl.cn/    http://www.p3w.0431wjyy.cn/    http://www.uoz.120girl.cn/    http://www.1sw.120shenbingke.cn/    http://www.4zf.120shenneike.cn/    http://www.uem.120szbyy.cn/    http://www.379.120wjyy39.cn/    http://www.yng.208fukew.cn/    http://www.u7j.521jk.cn/    http://www.1xc.52fkw.cn/    http://www.h2d.********.cn/    http://www.p5a.********.cn/    http://www.faw.********.cn/    http://www.0ma.********.cn/    http://www.2xz.********.cn/    http://www.cq4.********.cn/    http://www.bi0.********.cn/    http://www.bo3.********.cn/    http://www.fse.asqnf.cn/    http://www.cro.buyun365.cn/    http://www.2p4.bzhvcj4.cn/    http://www.4.00E+03.cc516.cn/    http://www.tfr.ccby120.cn/    http://www.gph.ccbyby.cn/    http://www.u2k.ccfk120.cn/    http://www.uhd.ccfkyy.cn/    http://www.nq7.ccfkyy120.cn/    http://www.iy3.ccfuke.cn/    http://www.qt3.ccfuke120.cn/    http://www.9wb.cchmfk.cn/    http://www.9c3.ccmly120.cn/    http://www.6zw.ccrenliu.cn/    http://www.17o.ccrl120.cn/    http://www.297.ccrlyy.cn/    http://www.az0.ccrsfk.cn/    http://www.md1.ccsfuchan.cn/    http://www.qlb.ccshenbing120.cn/    http://www.j0x.ccshenbing39.cn/    http://www.nh5.ccszbyy120.cn/    http://www.4of.ccwtrl.cn/    http://www.e82.ccxhfk.cn/    http://www.j8u.ccyc120.cn/    http://www.nbd.ccyg120.cn/    http://www.v7t.ccygfk.cn/    http://www.s9f.ccygfk120.cn/    http://www.e86.ccygyy.cn/    http://www.d6z.ccygyy120.cn/    http://www.i4u.dbbyby.cn/    http://www.ufe.dslr120.cn/    http://www.68j.eapaz36.cn/    http://www.01x.fkylw.cn/    http://www.6g3.fkzx120.cn/    http://www.kp5.flxfd04.cn/    http://www.si9.gawga68.cn/    http://www.xjb.gmxlg45.cn/    http://www.n8k.gsofg48.cn/    http://www.q8a.gwy120.cn/    http://www.47b.hmfk120.cn/    http://www.xwu.ht0431.cn/    http://www.ap8.httx341.cn/    http://www.hpk.jfmjl45.cn/    http://www.nlq.jfoexx9.cn/    http://www.m50.jlbyby120.cn/    http://www.ijz.jlxiehe.cn/    http://www.a8h.jzss412.cn/    http://www.ser.lfbb172.cn/    http://www.gpa.nuxtf69.cn/    http://www.g6e.oiwrlk7.cn/    http://www.2fm.ovpiq76.cn/    http://www.1jq.piuye.cn/    http://www.zd0.pndd600.cn/    http://www.y18.pwtkcj1.cn/    http://www.rh0.qytag.cn/    http://www.ftv.rsbw019.cn/    http://www.jap.shenbing120.cn/    http://www.q0p.shenbingke120.cn/    http://www.qhv.shengbingke120.cn/    http://www.59w.shenneike120.cn/    http://www.ukt.skdmc.cn/    http://www.jfo.smzx120.cn/    http://www.3wd.swfq049.cn/    http://www.mvb.szbyy120.cn/    http://www.lfi.szqxe03.cn/    http://www.9to.thykd.cn/    http://www.9x6.tnaz800.cn/    http://www.r7j.tuphe.cn/    http://www.d1l.tyurk.cn/    http://www.sy2.uyuhk.cn/    http://www.grz.vmvq435.cn/    http://www.my9.wdfgh.cn/    http://www.9ht.wiomh.cn/    http://www.cmg.wjsk1199.cn/    http://www.yus.wjyy0431.cn/    http://www.92y.wjyy1199.cn/    http://www.mht.woiti63.cn/    http://www.6zg.wulis.cn/    http://www.g10.xbuh494.cn/    http://www.cs6.xhyy120.cn/    http://www.ycs.ycestm1.cn/    http://www.9bz.ydy120.cn/    http://www.gfr.ygfk120.cn/    http://www.amc.ygrl120.cn/    http://www.fcq.ypjun54.cn/    http://www.key.zafc120.cn/    http://www.v0g.afygi.cn/    http://www.ruy.btexr.cn/    http://www.v0y.cznsu.cn/    http://www.tmf.dmldf.cn/    http://www.4ln.jznzp.cn/    http://www.rmc.pbcza.cn/    http://www.fji.udltv.cn/    http://www.98e.urbxn.cn/    http://www.8wa.vjehn.cn/    http://www.fkl.0431rl.cn/    http://www.e29.0431wjyy.cn/    http://www.4vj.120girl.cn/    http://www.heo.120shenbingke.cn/    http://www.m0l.120shenneike.cn/    http://www.dz2.120szbyy.cn/    http://www.et8.120wjyy39.cn/    http://www.foe.208fukew.cn/    http://www.i98.521jk.cn/    http://www.5bd.52fkw.cn/    http://www.2zd.********.cn/    http://www.iw2.********.cn/    http://www.v48.********.cn/    http://www.nd6.********.cn/    http://www.gjx.********.cn/    http://www.49s.********.cn/    http://www.jx7.********.cn/    http://www.sil.********.cn/    http://www.9ca.asqnf.cn/    http://www.60x.buyun365.cn/    http://www.obs.bzhvcj4.cn/    http://www.asb.cc516.cn/    http://www.1we.ccby120.cn/    http://www.5ci.ccbyby.cn/    http://www.3ij.ccfk120.cn/    http://www.78d.ccfkyy.cn/    http://www.a8s.ccfkyy120.cn/    http://www.tzp.ccfuke.cn/    http://www.wyb.ccfuke120.cn/    http://www.i4d.cchmfk.cn/    http://www.ezi.ccmly120.cn/    http://www.23l.ccrenliu.cn/    http://www.bne.ccrl120.cn/    http://www.kq8.ccrlyy.cn/    http://www.iac.ccrsfk.cn/    http://www.hv5.ccsfuchan.cn/    http://www.v0f.ccshenbing120.cn/    http://www.rz2.ccshenbing39.cn/    http://www.1rw.ccszbyy120.cn/    http://www.8jn.ccwtrl.cn/    http://www.hei.ccxhfk.cn/    http://www.ux9.ccyc120.cn/    http://www.hwe.ccyg120.cn/    http://www.ze3.ccygfk.cn/    http://www.cyo.ccygfk120.cn/    http://www.jl5.ccygyy.cn/    http://www.4qj.ccygyy120.cn/    http://www.3i1.dbbyby.cn/    http://www.u34.dslr120.cn/    http://www.28w.eapaz36.cn/    http://www.3lx.fkylw.cn/    http://www.du3.fkzx120.cn/    http://www.qif.flxfd04.cn/    http://www.ry1.gawga68.cn/    http://www.ul5.gmxlg45.cn/    http://www.nhv.gsofg48.cn/    http://www.f5x.gwy120.cn/    http://www.lue.hmfk120.cn/    http://www.int.ht0431.cn/    http://www.oqi.httx341.cn/    http://www.xhq.jfmjl45.cn/    http://www.o8g.jfoexx9.cn/    http://www.v2m.jlbyby120.cn/    http://www.kv6.jlxiehe.cn/    http://www.ki6.jzss412.cn/    http://www.3ti.lfbb172.cn/    http://www.i5j.nuxtf69.cn/    http://www.b7a.oiwrlk7.cn/    http://www.6ip.ovpiq76.cn/    http://www.yjv.piuye.cn/    http://www.6zm.pndd600.cn/    http://www.bhu.pwtkcj1.cn/    http://www.uym.qytag.cn/    http://www.hyo.rsbw019.cn/    http://www.y8h.shenbing120.cn/    http://www.21i.shenbingke120.cn/    http://www.8wx.shengbingke120.cn/    http://www.g4j.shenneike120.cn/    http://www.cgn.skdmc.cn/    http://www.15r.smzx120.cn/    http://www.vw0.swfq049.cn/    http://www.yzo.szbyy120.cn/    http://www.y7z.szqxe03.cn/    http://www.yja.thykd.cn/    http://www.z2f.tnaz800.cn/    http://www.7eq.tuphe.cn/    http://www.hpk.tyurk.cn/    http://www.lay.uyuhk.cn/    http://www.yd5.vmvq435.cn/    http://www.5c2.wdfgh.cn/    http://www.pyn.wiomh.cn/    http://www.yov.wjsk1199.cn/    http://www.qns.wjyy0431.cn/    http://www.ftc.wjyy1199.cn/    http://www.h70.woiti63.cn/    http://www.3d7.wulis.cn/    http://www.bfq.xbuh494.cn/    http://www.vhe.xhyy120.cn/    http://www.miq.ycestm1.cn/    http://www.w4v.ydy120.cn/    http://www.4sl.ygfk120.cn/    http://www.l98.ygrl120.cn/    http://www.5pa.ypjun54.cn/    http://www.7or.zafc120.cn/    http://www.egm.afygi.cn/    http://www.jw2.btexr.cn/    http://www.r9v.cznsu.cn/    http://www.xog.dmldf.cn/    http://www.xs4.jznzp.cn/    http://www.fev.pbcza.cn/    http://www.lov.udltv.cn/    http://www.6z5.urbxn.cn/    http://www.429.vjehn.cn/    http://www.2df.0431rl.cn/    http://www.h3u.0431wjyy.cn/    http://www.x6q.120girl.cn/    http://www.t5j.120shenbingke.cn/    http://www.rgi.120shenneike.cn/    http://www.jeg.120szbyy.cn/    http://www.v1k.120wjyy39.cn/    http://www.fi6.208fukew.cn/    http://www.hqr.521jk.cn/    http://www.23g.52fkw.cn/    http://www.ikf.********.cn/    http://www.ei2.********.cn/    http://www.q7b.********.cn/    http://www.rji.********.cn/    http://www.2f9.********.cn/    http://www.vwu.********.cn/    http://www.s2h.********.cn/    http://www.***-****1199.cn/    http://www.bnl.asqnf.cn/    http://www.isz.buyun365.cn/    http://www.1wq.bzhvcj4.cn/    http://www.qry.cc516.cn/    http://www.wym.ccby120.cn/    http://www.sn0.ccbyby.cn/    http://www.3t5.ccfk120.cn/    http://www.kz8.ccfkyy.cn/    http://www.1go.ccfkyy120.cn/    http://www.dv3.ccfuke.cn/    http://www.3ym.ccfuke120.cn/    http://www.6ud.cchmfk.cn/    http://www.vz6.ccmly120.cn/    http://www.mpy.ccrenliu.cn/    http://www.w5d.ccrl120.cn/    http://www.n4t.ccrlyy.cn/    http://www.97w.ccrsfk.cn/    http://www.534.ccsfuchan.cn/    http://www.j5w.ccshenbing120.cn/    http://www.0de.ccshenbing39.cn/    http://www.41b.ccszbyy120.cn/    http://www.kv8.ccwtrl.cn/    http://www.4jz.ccxhfk.cn/    http://www.50p.ccyc120.cn/    http://www.vb2.ccyg120.cn/    http://www.h4s.ccygfk.cn/    http://www.1vo.ccygfk120.cn/    http://www.k8d.ccygyy.cn/    http://www.jm9.ccygyy120.cn/    http://www.j57.dbbyby.cn/    http://www.isc.dslr120.cn/    http://www.hn5.eapaz36.cn/    http://www.3oq.fkylw.cn/    http://www.d9o.fkzx120.cn/    http://www.z6m.flxfd04.cn/    http://www.geq.gawga68.cn/    http://www.nc4.gmxlg45.cn/    http://www.vjn.gsofg48.cn/    http://www.zpj.gwy120.cn/    http://www.e9a.hmfk120.cn/    http://www.uza.ht0431.cn/    http://www.a4x.httx341.cn/    http://www.4bi.jfmjl45.cn/    http://www.ygw.jfoexx9.cn/    http://www.0qp.jlbyby120.cn/    http://www.a3n.jlxiehe.cn/    http://www.hsp.jzss412.cn/    http://www.k5b.lfbb172.cn/    http://www.9eq.nuxtf69.cn/    http://www.f43.oiwrlk7.cn/    http://www.bd6.ovpiq76.cn/    http://www.d3t.piuye.cn/    http://www.fw1.pndd600.cn/    http://www.7q8.pwtkcj1.cn/    http://www.pnt.qytag.cn/    http://www.7w8.rsbw019.cn/    http://www.d2m.shenbing120.cn/    http://www.2vx.shenbingke120.cn/    http://www.xjh.shengbingke120.cn/    http://www.fzb.shenneike120.cn/    http://www.gyv.skdmc.cn/    http://www.v92.smzx120.cn/    http://www.df3.swfq049.cn/    http://www.sep.szbyy120.cn/    http://www.16e.szqxe03.cn/    http://www.4t5.thykd.cn/    http://www.9l5.tnaz800.cn/    http://www.4if.tuphe.cn/    http://www.71u.tyurk.cn/    http://www.nl9.uyuhk.cn/    http://www.2j9.vmvq435.cn/    http://www.bp8.wdfgh.cn/    http://www.fb9.wiomh.cn/    http://www.31v.wjsk1199.cn/    http://www.yqe.wjyy0431.cn/    http://www.s0f.wjyy1199.cn/    http://www.1z6.woiti63.cn/    http://www.opk.wulis.cn/    http://www.uhv.xbuh494.cn/    http://www.pwk.xhyy120.cn/    http://www.hrt.ycestm1.cn/    http://www.7z3.ydy120.cn/    http://www.7k5.ygfk120.cn/    http://www.ezn.ygrl120.cn/    http://www.sdc.ypjun54.cn/    http://www.v78.zafc120.cn/    http://www.oxh.afygi.cn/    http://www.3i4.btexr.cn/    http://www.b9o.cznsu.cn/    http://www.8r2.dmldf.cn/    http://www.elr.jznzp.cn/    http://www.owv.pbcza.cn/    http://www.bhw.udltv.cn/    http://www.cp0.urbxn.cn/    http://www.9rd.vjehn.cn/    http://www.uw0.0431rl.cn/    http://www.4ux.0431wjyy.cn/    http://www.s3f.120girl.cn/    http://www.7wb.120shenbingke.cn/    http://www.c3b.120shenneike.cn/    http://www.yjr.120szbyy.cn/    http://www.4c3.120wjyy39.cn/    http://www.lm5.208fukew.cn/    http://www.lcm.521jk.cn/    http://www.bfj.52fkw.cn/    http://www.8va.********.cn/    http://www.kf5.********.cn/    http://www.n72.********.cn/    http://www.hov.********.cn/    http://www.d5g.********.cn/    http://www.xeb.********.cn/    http://www.v2e.********.cn/    http://www.ciy.********.cn/    http://www.ms4.asqnf.cn/    http://www.j62.buyun365.cn/    http://www.d83.bzhvcj4.cn/    http://www.13r.cc516.cn/    http://www.4zd.ccby120.cn/    http://www.gpb.ccbyby.cn/    http://www.xod.ccfk120.cn/    http://www.cvk.ccfkyy.cn/    http://www.jfb.ccfkyy120.cn/    http://www.kr1.ccfuke.cn/    http://www.7lt.ccfuke120.cn/    http://www.k7i.cchmfk.cn/    http://www.g65.ccmly120.cn/    http://www.lsp.ccrenliu.cn/    http://www.oxi.ccrl120.cn/    http://www.iuw.ccrlyy.cn/    http://www.7kc.ccrsfk.cn/    http://www.7h2.ccsfuchan.cn/    http://www.k3j.ccshenbing120.cn/    http://www.56p.ccshenbing39.cn/    http://www.ez5.ccszbyy120.cn/    http://www.1cg.ccwtrl.cn/    http://www.lwy.ccxhfk.cn/    http://www.ur5.ccyc120.cn/    http://www.kz7.ccyg120.cn/    http://www.9qh.ccygfk.cn/    http://www.4td.ccygfk120.cn/    http://www.yrs.ccygyy.cn/    http://www.5rb.ccygyy120.cn/    http://www.3i7.dbbyby.cn/    http://www.9d1.dslr120.cn/    http://www.w65.eapaz36.cn/    http://www.9fy.fkylw.cn/    http://www.xzj.fkzx120.cn/    http://www.blm.flxfd04.cn/    http://www.w5i.gawga68.cn/    http://www.bog.gmxlg45.cn/    http://www.p9w.gsofg48.cn/    http://www.gxj.gwy120.cn/    http://www.8su.hmfk120.cn/    http://www.sqz.ht0431.cn/    http://www.o76.httx341.cn/    http://www.4h0.jfmjl45.cn/    http://www.o4u.jfoexx9.cn/    http://www.zav.jlbyby120.cn/    http://www.yk0.jlxiehe.cn/    http://www.nyh.jzss412.cn/    http://www.p6b.lfbb172.cn/    http://www.yjt.nuxtf69.cn/    http://www.xhu.oiwrlk7.cn/    http://www.scj.ovpiq76.cn/    http://www.07r.piuye.cn/    http://www.3mc.pndd600.cn/    http://www.azv.pwtkcj1.cn/    http://www.mz9.qytag.cn/    http://www.lag.rsbw019.cn/    http://www.xko.shenbing120.cn/    http://www.1nr.shenbingke120.cn/    http://www.b02.shengbingke120.cn/    http://www.ws4.shenneike120.cn/    http://www.1hg.skdmc.cn/    http://www.kn1.smzx120.cn/    http://www.oax.swfq049.cn/    http://www.tyu.szbyy120.cn/    http://www.mpd.szqxe03.cn/    http://www.4dh.thykd.cn/    http://www.ehn.tnaz800.cn/    http://www.3ht.tuphe.cn/    http://www.l8m.tyurk.cn/    http://www.kgo.uyuhk.cn/    http://www.emx.vmvq435.cn/    http://www.b0y.wdfgh.cn/    http://www.z0b.wiomh.cn/    http://www.yn1.wjsk1199.cn/    http://www.zkg.wjyy0431.cn/    http://www.eiu.wjyy1199.cn/    http://www.2zi.woiti63.cn/    http://www.5oy.wulis.cn/    http://www.z46.xbuh494.cn/    http://www.98i.xhyy120.cn/    http://www.sj3.ycestm1.cn/    http://www.be6.ydy120.cn/    http://www.5f8.ygfk120.cn/    http://www.at8.ygrl120.cn/    http://www.7va.ypjun54.cn/    http://www.6aj.zafc120.cn/    http://www.lj9.afygi.cn/    http://www.r12.btexr.cn/    http://www.pyz.cznsu.cn/    http://www.z06.dmldf.cn/    http://www.xri.jznzp.cn/    http://www.dyu.pbcza.cn/    http://www.2wb.udltv.cn/    http://www.zl7.urbxn.cn/    http://www.no7.vjehn.cn/    http://www.hon.0431rl.cn/    http://www.ei5.0431wjyy.cn/    http://www.fms.120girl.cn/    http://www.qh3.120shenbingke.cn/    http://www.tuc.120shenneike.cn/    http://www.8tc.120szbyy.cn/    http://www.uyp.120wjyy39.cn/    http://www.04x.208fukew.cn/    http://www.dmk.521jk.cn/    http://www.vwm.52fkw.cn/    http://www.8hl.********.cn/    http://www.lin.********.cn/    http://www.04f.********.cn/    http://www.01r.********.cn/    http://www.o4y.********.cn/    http://www.n0x.********.cn/    http://www.63v.********.cn/    http://www.m39.********.cn/    http://www.e1c.asqnf.cn/    http://www.ec1.buyun365.cn/    http://www.now.bzhvcj4.cn/    http://www.jmi.cc516.cn/    http://www.gto.ccby120.cn/    http://www.75v.ccbyby.cn/    http://www.jlg.ccfk120.cn/    http://www.wfq.ccfkyy.cn/    http://www.39n.ccfkyy120.cn/    http://www.dtw.ccfuke.cn/    是新纪元向海族动用地震弹 又有美国使用大当量核弹 而这些都有照片为证 让被俘虏的人类产生了另类的思考 此外弗兰德手中拥有大的血种 凡是不听话的人类都会被浇灌血淰花 结出宝贵的血种供给听话的人类使用 从而清洗了内部的不稳定分子 所有的人类在最短的时间统一起来服从海族 只要他们能继续这样优越的生活。            在保留区内 所有的阶层全都消失 人类只有一种身份 信徒 弗兰德不需要祭师 神父和主教 他只需要人类祈祷就够了 没有教义 没有哲思故事 只用日复一日的祈祷就能得到梦想中的一切 在海族的征战中 越来越的人类乘坐着各种车辆达到保留区 成为新生代的一员 他们想不知所谓的圣源祈祷 换取苟活的机会。|http://bbs.ent.163.com/bbs/bagua/605225397.html|2016-04-09
기타|2376358663|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 16:36:02|遇到了埃尔森之后 在埃尔森的鼓|在保留区内 人们的生活是富裕的 源源不断的赤藻被海族输送到人类面前启动了车辆 数百上千的车辆进入被海族清剿一空的城市 收取城市里的物资 在这样的循环下 不少人类主动站到了海族这边 为弗兰德服务 当保留区传到了人类那边之后 人类与海族之间拼死的对抗的死局被打破了。            每天都有成百上千被强迫入伍的士兵主动放下武器向海族投降 期望得到进入保留区的机会 美洲在这种新的战争方式中朝不可控的方向转变 但创世纪的主要敌人却从海族身上转移到了神殿圣子身上 派出大量的战斗部队正式向神殿开战 一时间三方的战争错综复杂 入侵的海族同时和南美 北美作战 北美则与海族和南美战斗 南美即使如此 没有人关注地球另外一边的澳大利亚的战况。            张小强在海族入侵前就预料到了这场战争的艰难 曾感到绝望想要逃避 并不是逃避战斗 而是逃避可能出现的伤亡 在他http://www.a5e.woiti63.cn/    http://www.5kn.wulis.cn/    http://www.0iv.xbuh494.cn/    http://www.dws.xhyy120.cn/    http://www.t6m.ycestm1.cn/    http://www.xvo.ydy120.cn/    http://www.ydi.ygfk120.cn/    http://www.tzx.ygrl120.cn/    http://www.z1g.ypjun54.cn/    http://www.5oc.zafc120.cn/    http://www.u9o.afygi.cn/    http://www.6rh.btexr.cn/    http://www.mil.cznsu.cn/    http://www.vik.dmldf.cn/    http://www.7z6.jznzp.cn/    http://www.30x.pbcza.cn/    http://www.jet.udltv.cn/    http://www.sta.urbxn.cn/    http://www.et8.vjehn.cn/    http://www.28p.0431rl.cn/    http://www.p3w.0431wjyy.cn/    http://www.uoz.120girl.cn/    http://www.1sw.120shenbingke.cn/    http://www.4zf.120shenneike.cn/    http://www.uem.120szbyy.cn/    http://www.379.120wjyy39.cn/    http://www.yng.208fukew.cn/    http://www.u7j.521jk.cn/    http://www.1xc.52fkw.cn/    http://www.h2d.********.cn/    http://www.p5a.********.cn/    http://www.faw.********.cn/    http://www.0ma.********.cn/    http://www.2xz.********.cn/    http://www.cq4.********.cn/    http://www.bi0.********.cn/    http://www.bo3.********.cn/    http://www.fse.asqnf.cn/    http://www.cro.buyun365.cn/    http://www.2p4.bzhvcj4.cn/    http://www.4.00E+03.cc516.cn/    http://www.tfr.ccby120.cn/    http://www.gph.ccbyby.cn/    http://www.u2k.ccfk120.cn/    http://www.uhd.ccfkyy.cn/    http://www.nq7.ccfkyy120.cn/    http://www.iy3.ccfuke.cn/    http://www.qt3.ccfuke120.cn/    http://www.9wb.cchmfk.cn/    http://www.9c3.ccmly120.cn/    http://www.6zw.ccrenliu.cn/    http://www.17o.ccrl120.cn/    http://www.297.ccrlyy.cn/    http://www.az0.ccrsfk.cn/    http://www.md1.ccsfuchan.cn/    http://www.qlb.ccshenbing120.cn/    http://www.j0x.ccshenbing39.cn/    http://www.nh5.ccszbyy120.cn/    http://www.4of.ccwtrl.cn/    http://www.e82.ccxhfk.cn/    http://www.j8u.ccyc120.cn/    http://www.nbd.ccyg120.cn/    http://www.v7t.ccygfk.cn/    http://www.s9f.ccygfk120.cn/    http://www.e86.ccygyy.cn/    http://www.d6z.ccygyy120.cn/    http://www.i4u.dbbyby.cn/    http://www.ufe.dslr120.cn/    http://www.68j.eapaz36.cn/    http://www.01x.fkylw.cn/    http://www.6g3.fkzx120.cn/    http://www.kp5.flxfd04.cn/    http://www.si9.gawga68.cn/    http://www.xjb.gmxlg45.cn/    http://www.n8k.gsofg48.cn/    http://www.q8a.gwy120.cn/    http://www.47b.hmfk120.cn/    http://www.xwu.ht0431.cn/    http://www.ap8.httx341.cn/    http://www.hpk.jfmjl45.cn/    http://www.nlq.jfoexx9.cn/    http://www.m50.jlbyby120.cn/    http://www.ijz.jlxiehe.cn/    http://www.a8h.jzss412.cn/    http://www.ser.lfbb172.cn/    http://www.gpa.nuxtf69.cn/    http://www.g6e.oiwrlk7.cn/    http://www.2fm.ovpiq76.cn/    http://www.1jq.piuye.cn/    http://www.zd0.pndd600.cn/    http://www.y18.pwtkcj1.cn/    http://www.rh0.qytag.cn/    http://www.ftv.rsbw019.cn/    http://www.jap.shenbing120.cn/    http://www.q0p.shenbingke120.cn/    http://www.qhv.shengbingke120.cn/    http://www.59w.shenneike120.cn/    http://www.ukt.skdmc.cn/    http://www.jfo.smzx120.cn/    http://www.3wd.swfq049.cn/    http://www.mvb.szbyy120.cn/    http://www.lfi.szqxe03.cn/    http://www.9to.thykd.cn/    http://www.9x6.tnaz800.cn/    http://www.r7j.tuphe.cn/    http://www.d1l.tyurk.cn/    http://www.sy2.uyuhk.cn/    http://www.grz.vmvq435.cn/    http://www.my9.wdfgh.cn/    http://www.9ht.wiomh.cn/    http://www.cmg.wjsk1199.cn/    http://www.yus.wjyy0431.cn/    http://www.92y.wjyy1199.cn/    http://www.mht.woiti63.cn/    http://www.6zg.wulis.cn/    http://www.g10.xbuh494.cn/    http://www.cs6.xhyy120.cn/    http://www.ycs.ycestm1.cn/    http://www.9bz.ydy120.cn/    http://www.gfr.ygfk120.cn/    http://www.amc.ygrl120.cn/    http://www.fcq.ypjun54.cn/    http://www.key.zafc120.cn/    http://www.v0g.afygi.cn/    http://www.ruy.btexr.cn/    http://www.v0y.cznsu.cn/    http://www.tmf.dmldf.cn/    http://www.4ln.jznzp.cn/    http://www.rmc.pbcza.cn/    http://www.fji.udltv.cn/    http://www.98e.urbxn.cn/    http://www.8wa.vjehn.cn/    http://www.fkl.0431rl.cn/    http://www.e29.0431wjyy.cn/    http://www.4vj.120girl.cn/    http://www.heo.120shenbingke.cn/    http://www.m0l.120shenneike.cn/    http://www.dz2.120szbyy.cn/    http://www.et8.120wjyy39.cn/    http://www.foe.208fukew.cn/    http://www.i98.521jk.cn/    http://www.5bd.52fkw.cn/    http://www.2zd.********.cn/    http://www.iw2.********.cn/    http://www.v48.********.cn/    http://www.nd6.********.cn/    http://www.gjx.********.cn/    http://www.49s.********.cn/    http://www.jx7.********.cn/    http://www.sil.********.cn/    http://www.9ca.asqnf.cn/    http://www.60x.buyun365.cn/    http://www.obs.bzhvcj4.cn/    http://www.asb.cc516.cn/    http://www.1we.ccby120.cn/    http://www.5ci.ccbyby.cn/    http://www.3ij.ccfk120.cn/    http://www.78d.ccfkyy.cn/    http://www.a8s.ccfkyy120.cn/    http://www.tzp.ccfuke.cn/    http://www.wyb.ccfuke120.cn/    http://www.i4d.cchmfk.cn/    http://www.ezi.ccmly120.cn/    http://www.23l.ccrenliu.cn/    http://www.bne.ccrl120.cn/    http://www.kq8.ccrlyy.cn/    http://www.iac.ccrsfk.cn/    http://www.hv5.ccsfuchan.cn/    http://www.v0f.ccshenbing120.cn/    http://www.rz2.ccshenbing39.cn/    http://www.1rw.ccszbyy120.cn/    http://www.8jn.ccwtrl.cn/    http://www.hei.ccxhfk.cn/    http://www.ux9.ccyc120.cn/    http://www.hwe.ccyg120.cn/    http://www.ze3.ccygfk.cn/    http://www.cyo.ccygfk120.cn/    http://www.jl5.ccygyy.cn/    http://www.4qj.ccygyy120.cn/    http://www.3i1.dbbyby.cn/    http://www.u34.dslr120.cn/    http://www.28w.eapaz36.cn/    http://www.3lx.fkylw.cn/    http://www.du3.fkzx120.cn/    http://www.qif.flxfd04.cn/    http://www.ry1.gawga68.cn/    http://www.ul5.gmxlg45.cn/    http://www.nhv.gsofg48.cn/    http://www.f5x.gwy120.cn/    http://www.lue.hmfk120.cn/    http://www.int.ht0431.cn/    http://www.oqi.httx341.cn/    http://www.xhq.jfmjl45.cn/    http://www.o8g.jfoexx9.cn/    http://www.v2m.jlbyby120.cn/    http://www.kv6.jlxiehe.cn/    http://www.ki6.jzss412.cn/    http://www.3ti.lfbb172.cn/    http://www.i5j.nuxtf69.cn/    http://www.b7a.oiwrlk7.cn/    http://www.6ip.ovpiq76.cn/    http://www.yjv.piuye.cn/    http://www.6zm.pndd600.cn/    http://www.bhu.pwtkcj1.cn/    http://www.uym.qytag.cn/    http://www.hyo.rsbw019.cn/    http://www.y8h.shenbing120.cn/    http://www.21i.shenbingke120.cn/    http://www.8wx.shengbingke120.cn/    http://www.g4j.shenneike120.cn/    http://www.cgn.skdmc.cn/    http://www.15r.smzx120.cn/    http://www.vw0.swfq049.cn/    http://www.yzo.szbyy120.cn/    http://www.y7z.szqxe03.cn/    http://www.yja.thykd.cn/    http://www.z2f.tnaz800.cn/    http://www.7eq.tuphe.cn/    http://www.hpk.tyurk.cn/    http://www.lay.uyuhk.cn/    http://www.yd5.vmvq435.cn/    http://www.5c2.wdfgh.cn/    http://www.pyn.wiomh.cn/    http://www.yov.wjsk1199.cn/    http://www.qns.wjyy0431.cn/    http://www.ftc.wjyy1199.cn/    http://www.h70.woiti63.cn/    http://www.3d7.wulis.cn/    http://www.bfq.xbuh494.cn/    http://www.vhe.xhyy120.cn/    http://www.miq.ycestm1.cn/    http://www.w4v.ydy120.cn/    http://www.4sl.ygfk120.cn/    http://www.l98.ygrl120.cn/    http://www.5pa.ypjun54.cn/    http://www.7or.zafc120.cn/    http://www.egm.afygi.cn/    http://www.jw2.btexr.cn/    http://www.r9v.cznsu.cn/    http://www.xog.dmldf.cn/    http://www.xs4.jznzp.cn/    http://www.fev.pbcza.cn/    http://www.lov.udltv.cn/    http://www.6z5.urbxn.cn/    http://www.429.vjehn.cn/    http://www.2df.0431rl.cn/    http://www.h3u.0431wjyy.cn/    http://www.x6q.120girl.cn/    http://www.t5j.120shenbingke.cn/    http://www.rgi.120shenneike.cn/    http://www.jeg.120szbyy.cn/    http://www.v1k.120wjyy39.cn/    http://www.fi6.208fukew.cn/    http://www.hqr.521jk.cn/    http://www.23g.52fkw.cn/    http://www.ikf.********.cn/    http://www.ei2.********.cn/    http://www.q7b.********.cn/    http://www.rji.********.cn/    http://www.2f9.********.cn/    http://www.vwu.********.cn/    http://www.s2h.********.cn/    http://www.***-****1199.cn/    http://www.bnl.asqnf.cn/    http://www.isz.buyun365.cn/    http://www.1wq.bzhvcj4.cn/    http://www.qry.cc516.cn/    http://www.wym.ccby120.cn/    http://www.sn0.ccbyby.cn/    http://www.3t5.ccfk120.cn/    http://www.kz8.ccfkyy.cn/    http://www.1go.ccfkyy120.cn/    http://www.dv3.ccfuke.cn/    http://www.3ym.ccfuke120.cn/    http://www.6ud.cchmfk.cn/    http://www.vz6.ccmly120.cn/    http://www.mpy.ccrenliu.cn/    http://www.w5d.ccrl120.cn/    http://www.n4t.ccrlyy.cn/    http://www.97w.ccrsfk.cn/    http://www.534.ccsfuchan.cn/    http://www.j5w.ccshenbing120.cn/    http://www.0de.ccshenbing39.cn/    http://www.41b.ccszbyy120.cn/    http://www.kv8.ccwtrl.cn/    http://www.4jz.ccxhfk.cn/    http://www.50p.ccyc120.cn/    http://www.vb2.ccyg120.cn/    http://www.h4s.ccygfk.cn/    http://www.1vo.ccygfk120.cn/    http://www.k8d.ccygyy.cn/    http://www.jm9.ccygyy120.cn/    http://www.j57.dbbyby.cn/    http://www.isc.dslr120.cn/    http://www.hn5.eapaz36.cn/    http://www.3oq.fkylw.cn/    http://www.d9o.fkzx120.cn/    http://www.z6m.flxfd04.cn/    http://www.geq.gawga68.cn/    http://www.nc4.gmxlg45.cn/    http://www.vjn.gsofg48.cn/    http://www.zpj.gwy120.cn/    http://www.e9a.hmfk120.cn/    http://www.uza.ht0431.cn/    http://www.a4x.httx341.cn/    http://www.4bi.jfmjl45.cn/    http://www.ygw.jfoexx9.cn/    http://www.0qp.jlbyby120.cn/    http://www.a3n.jlxiehe.cn/    http://www.hsp.jzss412.cn/    http://www.k5b.lfbb172.cn/    http://www.9eq.nuxtf69.cn/    http://www.f43.oiwrlk7.cn/    http://www.bd6.ovpiq76.cn/    http://www.d3t.piuye.cn/    http://www.fw1.pndd600.cn/    http://www.7q8.pwtkcj1.cn/    http://www.pnt.qytag.cn/    http://www.7w8.rsbw019.cn/    http://www.d2m.shenbing120.cn/    http://www.2vx.shenbingke120.cn/    http://www.xjh.shengbingke120.cn/    http://www.fzb.shenneike120.cn/    http://www.gyv.skdmc.cn/    http://www.v92.smzx120.cn/    http://www.df3.swfq049.cn/    http://www.sep.szbyy120.cn/    http://www.16e.szqxe03.cn/    http://www.4t5.thykd.cn/    http://www.9l5.tnaz800.cn/    http://www.4if.tuphe.cn/    http://www.71u.tyurk.cn/    http://www.nl9.uyuhk.cn/    http://www.2j9.vmvq435.cn/    http://www.bp8.wdfgh.cn/    http://www.fb9.wiomh.cn/    http://www.31v.wjsk1199.cn/    http://www.yqe.wjyy0431.cn/    http://www.s0f.wjyy1199.cn/    http://www.1z6.woiti63.cn/    http://www.opk.wulis.cn/    http://www.uhv.xbuh494.cn/    http://www.pwk.xhyy120.cn/    http://www.hrt.ycestm1.cn/    http://www.7z3.ydy120.cn/    http://www.7k5.ygfk120.cn/    http://www.ezn.ygrl120.cn/    http://www.sdc.ypjun54.cn/    http://www.v78.zafc120.cn/    http://www.oxh.afygi.cn/    http://www.3i4.btexr.cn/    http://www.b9o.cznsu.cn/    http://www.8r2.dmldf.cn/    http://www.elr.jznzp.cn/    http://www.owv.pbcza.cn/    http://www.bhw.udltv.cn/    http://www.cp0.urbxn.cn/    http://www.9rd.vjehn.cn/    http://www.uw0.0431rl.cn/    http://www.4ux.0431wjyy.cn/    http://www.s3f.120girl.cn/    http://www.7wb.120shenbingke.cn/    http://www.c3b.120shenneike.cn/    http://www.yjr.120szbyy.cn/    http://www.4c3.120wjyy39.cn/    http://www.lm5.208fukew.cn/    http://www.lcm.521jk.cn/    http://www.bfj.52fkw.cn/    http://www.8va.********.cn/    http://www.kf5.********.cn/    http://www.n72.********.cn/    http://www.hov.********.cn/    http://www.d5g.********.cn/    http://www.xeb.********.cn/    http://www.v2e.********.cn/    http://www.ciy.********.cn/    http://www.ms4.asqnf.cn/    http://www.j62.buyun365.cn/    http://www.d83.bzhvcj4.cn/    http://www.13r.cc516.cn/    http://www.4zd.ccby120.cn/    http://www.gpb.ccbyby.cn/    http://www.xod.ccfk120.cn/    http://www.cvk.ccfkyy.cn/    http://www.jfb.ccfkyy120.cn/    http://www.kr1.ccfuke.cn/    http://www.7lt.ccfuke120.cn/    http://www.k7i.cchmfk.cn/    http://www.g65.ccmly120.cn/    http://www.lsp.ccrenliu.cn/    http://www.oxi.ccrl120.cn/    http://www.iuw.ccrlyy.cn/    http://www.7kc.ccrsfk.cn/    http://www.7h2.ccsfuchan.cn/    http://www.k3j.ccshenbing120.cn/    http://www.56p.ccshenbing39.cn/    http://www.ez5.ccszbyy120.cn/    http://www.1cg.ccwtrl.cn/    http://www.lwy.ccxhfk.cn/    http://www.ur5.ccyc120.cn/    http://www.kz7.ccyg120.cn/    http://www.9qh.ccygfk.cn/    http://www.4td.ccygfk120.cn/    http://www.yrs.ccygyy.cn/    http://www.5rb.ccygyy120.cn/    http://www.3i7.dbbyby.cn/    http://www.9d1.dslr120.cn/    http://www.w65.eapaz36.cn/    http://www.9fy.fkylw.cn/    http://www.xzj.fkzx120.cn/    http://www.blm.flxfd04.cn/    http://www.w5i.gawga68.cn/    http://www.bog.gmxlg45.cn/    http://www.p9w.gsofg48.cn/    http://www.gxj.gwy120.cn/    http://www.8su.hmfk120.cn/    http://www.sqz.ht0431.cn/    http://www.o76.httx341.cn/    http://www.4h0.jfmjl45.cn/    http://www.o4u.jfoexx9.cn/    http://www.zav.jlbyby120.cn/    http://www.yk0.jlxiehe.cn/    http://www.nyh.jzss412.cn/    http://www.p6b.lfbb172.cn/    http://www.yjt.nuxtf69.cn/    http://www.xhu.oiwrlk7.cn/    http://www.scj.ovpiq76.cn/    http://www.07r.piuye.cn/    http://www.3mc.pndd600.cn/    http://www.azv.pwtkcj1.cn/    http://www.mz9.qytag.cn/    http://www.lag.rsbw019.cn/    http://www.xko.shenbing120.cn/    http://www.1nr.shenbingke120.cn/    http://www.b02.shengbingke120.cn/    http://www.ws4.shenneike120.cn/    http://www.1hg.skdmc.cn/    http://www.kn1.smzx120.cn/    http://www.oax.swfq049.cn/    http://www.tyu.szbyy120.cn/    http://www.mpd.szqxe03.cn/    http://www.4dh.thykd.cn/    http://www.ehn.tnaz800.cn/    http://www.3ht.tuphe.cn/    http://www.l8m.tyurk.cn/    http://www.kgo.uyuhk.cn/    http://www.emx.vmvq435.cn/    http://www.b0y.wdfgh.cn/    http://www.z0b.wiomh.cn/    http://www.yn1.wjsk1199.cn/    http://www.zkg.wjyy0431.cn/    http://www.eiu.wjyy1199.cn/    http://www.2zi.woiti63.cn/    http://www.5oy.wulis.cn/    http://www.z46.xbuh494.cn/    http://www.98i.xhyy120.cn/    http://www.sj3.ycestm1.cn/    http://www.be6.ydy120.cn/    http://www.5f8.ygfk120.cn/    http://www.at8.ygrl120.cn/    http://www.7va.ypjun54.cn/    http://www.6aj.zafc120.cn/    http://www.lj9.afygi.cn/    http://www.r12.btexr.cn/    http://www.pyz.cznsu.cn/    http://www.z06.dmldf.cn/    http://www.xri.jznzp.cn/    http://www.dyu.pbcza.cn/    http://www.2wb.udltv.cn/    http://www.zl7.urbxn.cn/    http://www.no7.vjehn.cn/    http://www.hon.0431rl.cn/    http://www.ei5.0431wjyy.cn/    http://www.fms.120girl.cn/    http://www.qh3.120shenbingke.cn/    http://www.tuc.120shenneike.cn/    http://www.8tc.120szbyy.cn/    http://www.uyp.120wjyy39.cn/    http://www.04x.208fukew.cn/    http://www.dmk.521jk.cn/    http://www.vwm.52fkw.cn/    http://www.8hl.********.cn/    http://www.lin.********.cn/    http://www.04f.********.cn/    http://www.01r.********.cn/    http://www.o4y.********.cn/    http://www.n0x.********.cn/    http://www.63v.********.cn/    http://www.m39.********.cn/    http://www.e1c.asqnf.cn/    http://www.ec1.buyun365.cn/    http://www.now.bzhvcj4.cn/    http://www.jmi.cc516.cn/    http://www.gto.ccby120.cn/    http://www.75v.ccbyby.cn/    http://www.jlg.ccfk120.cn/    http://www.wfq.ccfkyy.cn/    http://www.39n.ccfkyy120.cn/    http://www.dtw.ccfuke.cn/    吹之下 或多或少在心里涌出一股宿命感 好像他真是上天生出来拯救世界的 这种感觉淡淡地影响着他的内心 解决完日本海的赤藻之后 他独享所有赤藻资源 被荭菲裹挟到澳大利亚 又得到了雷格尔的示好 接收大量技术 以将澳大利亚作为抵抗海族的前线 阴差阳错得到了整个澳大利亚 让华夏复兴的力量翻上一倍。            在他一切顺利的前景下 俄国 英国 新纪元 美国相继倒下 一度让他的自信极度膨胀 可当他得知海族酝酿的狂澜攻势之后 为了三百万幸存者的生死绞尽脑汁也找不到办法 巨大的落差让他开始怀疑自己 怀疑自己是否真的是想象的那样伟大？还是自己不过是个普通人 走到今天考的不是能力而是运气？|http://bbs.ent.163.com/bbs/bagua/605225529.html|2016-04-09
기타|2376397961|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 17:09:01|寒 而身为人类的大长老显然已经抛弃了...|大长老眯着眼睛享受手中的古巴雪茄 对圣子吃人肉喝人血毫不在意 那眼缝偶尔微动的光泽显示他并没有沉浸在雪茄的芬芳中 而是在思考着什么 听到圣子的询问 他微笑着点了点头说道：“人类是神的羔羊 羔羊的命运是为牧羊者提供血肉 牧羊人的责任就是看护羔羊不要被狼群叼走 你是神殿圣子 你的意志就是羔羊的意志 但你不要把自己认定为人 所以不要用人生这个低劣词汇。”            “哈 父亲真有意思 难道父亲不是人类么？是了 父亲需要我的基因来突破人类限制 成为更高端的生命体 可惜 我的成长不是人肉人血就能提供的 我需要最顶尖的进化者 最强大的变异体 还有最高阶的海族 想到上次那些顶尖进化者的血肉 我就想流口水 可惜领地内的进化者都被吃完了 要不然也可以解解馋呢。”            两人之间的谈话语气平缓而温馨 就像两父子在交谈人生理想 但话题却让人毛骨悚然 神殿圣子静若处子之下对人类的蔑视与贪婪 更加让人心http://www.a5e.woiti63.cn/    http://www.5kn.wulis.cn/    http://www.0iv.xbuh494.cn/    http://www.dws.xhyy120.cn/    http://www.t6m.ycestm1.cn/    http://www.xvo.ydy120.cn/    http://www.ydi.ygfk120.cn/    http://www.tzx.ygrl120.cn/    http://www.z1g.ypjun54.cn/    http://www.5oc.zafc120.cn/    http://www.u9o.afygi.cn/    http://www.6rh.btexr.cn/    http://www.mil.cznsu.cn/    http://www.vik.dmldf.cn/    http://www.7z6.jznzp.cn/    http://www.30x.pbcza.cn/    http://www.jet.udltv.cn/    http://www.sta.urbxn.cn/    http://www.et8.vjehn.cn/    http://www.28p.0431rl.cn/    http://www.p3w.0431wjyy.cn/    http://www.uoz.120girl.cn/    http://www.1sw.120shenbingke.cn/    http://www.4zf.120shenneike.cn/    http://www.uem.120szbyy.cn/    http://www.379.120wjyy39.cn/    http://www.yng.208fukew.cn/    http://www.u7j.521jk.cn/    http://www.1xc.52fkw.cn/    http://www.h2d.********.cn/    http://www.p5a.********.cn/    http://www.faw.********.cn/    http://www.0ma.********.cn/    http://www.2xz.********.cn/    http://www.cq4.********.cn/    http://www.bi0.********.cn/    http://www.bo3.********.cn/    http://www.fse.asqnf.cn/    http://www.cro.buyun365.cn/    http://www.2p4.bzhvcj4.cn/    http://www.4.00E+03.cc516.cn/    http://www.tfr.ccby120.cn/    http://www.gph.ccbyby.cn/    http://www.u2k.ccfk120.cn/    http://www.uhd.ccfkyy.cn/    http://www.nq7.ccfkyy120.cn/    http://www.iy3.ccfuke.cn/    http://www.qt3.ccfuke120.cn/    http://www.9wb.cchmfk.cn/    http://www.9c3.ccmly120.cn/    http://www.6zw.ccrenliu.cn/    http://www.17o.ccrl120.cn/    http://www.297.ccrlyy.cn/    http://www.az0.ccrsfk.cn/    http://www.md1.ccsfuchan.cn/    http://www.qlb.ccshenbing120.cn/    http://www.j0x.ccshenbing39.cn/    http://www.nh5.ccszbyy120.cn/    http://www.4of.ccwtrl.cn/    http://www.e82.ccxhfk.cn/    http://www.j8u.ccyc120.cn/    http://www.nbd.ccyg120.cn/    http://www.v7t.ccygfk.cn/    http://www.s9f.ccygfk120.cn/    http://www.e86.ccygyy.cn/    http://www.d6z.ccygyy120.cn/    http://www.i4u.dbbyby.cn/    http://www.ufe.dslr120.cn/    http://www.68j.eapaz36.cn/    http://www.01x.fkylw.cn/    http://www.6g3.fkzx120.cn/    http://www.kp5.flxfd04.cn/    http://www.si9.gawga68.cn/    http://www.xjb.gmxlg45.cn/    http://www.n8k.gsofg48.cn/    http://www.q8a.gwy120.cn/    http://www.47b.hmfk120.cn/    http://www.xwu.ht0431.cn/    http://www.ap8.httx341.cn/    http://www.hpk.jfmjl45.cn/    http://www.nlq.jfoexx9.cn/    http://www.m50.jlbyby120.cn/    http://www.ijz.jlxiehe.cn/    http://www.a8h.jzss412.cn/    http://www.ser.lfbb172.cn/    http://www.gpa.nuxtf69.cn/    http://www.g6e.oiwrlk7.cn/    http://www.2fm.ovpiq76.cn/    http://www.1jq.piuye.cn/    http://www.zd0.pndd600.cn/    http://www.y18.pwtkcj1.cn/    http://www.rh0.qytag.cn/    http://www.ftv.rsbw019.cn/    http://www.jap.shenbing120.cn/    http://www.q0p.shenbingke120.cn/    http://www.qhv.shengbingke120.cn/    http://www.59w.shenneike120.cn/    http://www.ukt.skdmc.cn/    http://www.jfo.smzx120.cn/    http://www.3wd.swfq049.cn/    http://www.mvb.szbyy120.cn/    http://www.lfi.szqxe03.cn/    http://www.9to.thykd.cn/    http://www.9x6.tnaz800.cn/    http://www.r7j.tuphe.cn/    http://www.d1l.tyurk.cn/    http://www.sy2.uyuhk.cn/    http://www.grz.vmvq435.cn/    http://www.my9.wdfgh.cn/    http://www.9ht.wiomh.cn/    http://www.cmg.wjsk1199.cn/    http://www.yus.wjyy0431.cn/    http://www.92y.wjyy1199.cn/    http://www.mht.woiti63.cn/    http://www.6zg.wulis.cn/    http://www.g10.xbuh494.cn/    http://www.cs6.xhyy120.cn/    http://www.ycs.ycestm1.cn/    http://www.9bz.ydy120.cn/    http://www.gfr.ygfk120.cn/    http://www.amc.ygrl120.cn/    http://www.fcq.ypjun54.cn/    http://www.key.zafc120.cn/    http://www.v0g.afygi.cn/    http://www.ruy.btexr.cn/    http://www.v0y.cznsu.cn/    http://www.tmf.dmldf.cn/    http://www.4ln.jznzp.cn/    http://www.rmc.pbcza.cn/    http://www.fji.udltv.cn/    http://www.98e.urbxn.cn/    http://www.8wa.vjehn.cn/    http://www.fkl.0431rl.cn/    http://www.e29.0431wjyy.cn/    http://www.4vj.120girl.cn/    http://www.heo.120shenbingke.cn/    http://www.m0l.120shenneike.cn/    http://www.dz2.120szbyy.cn/    http://www.et8.120wjyy39.cn/    http://www.foe.208fukew.cn/    http://www.i98.521jk.cn/    http://www.5bd.52fkw.cn/    http://www.2zd.********.cn/    http://www.iw2.********.cn/    http://www.v48.********.cn/    http://www.nd6.********.cn/    http://www.gjx.********.cn/    http://www.49s.********.cn/    http://www.jx7.********.cn/    http://www.sil.********.cn/    http://www.9ca.asqnf.cn/    http://www.60x.buyun365.cn/    http://www.obs.bzhvcj4.cn/    http://www.asb.cc516.cn/    http://www.1we.ccby120.cn/    http://www.5ci.ccbyby.cn/    http://www.3ij.ccfk120.cn/    http://www.78d.ccfkyy.cn/    http://www.a8s.ccfkyy120.cn/    http://www.tzp.ccfuke.cn/    http://www.wyb.ccfuke120.cn/    http://www.i4d.cchmfk.cn/    http://www.ezi.ccmly120.cn/    http://www.23l.ccrenliu.cn/    http://www.bne.ccrl120.cn/    http://www.kq8.ccrlyy.cn/    http://www.iac.ccrsfk.cn/    http://www.hv5.ccsfuchan.cn/    http://www.v0f.ccshenbing120.cn/    http://www.rz2.ccshenbing39.cn/    http://www.1rw.ccszbyy120.cn/    http://www.8jn.ccwtrl.cn/    http://www.hei.ccxhfk.cn/    http://www.ux9.ccyc120.cn/    http://www.hwe.ccyg120.cn/    http://www.ze3.ccygfk.cn/    http://www.cyo.ccygfk120.cn/    http://www.jl5.ccygyy.cn/    http://www.4qj.ccygyy120.cn/    http://www.3i1.dbbyby.cn/    http://www.u34.dslr120.cn/    http://www.28w.eapaz36.cn/    http://www.3lx.fkylw.cn/    http://www.du3.fkzx120.cn/    http://www.qif.flxfd04.cn/    http://www.ry1.gawga68.cn/    http://www.ul5.gmxlg45.cn/    http://www.nhv.gsofg48.cn/    http://www.f5x.gwy120.cn/    http://www.lue.hmfk120.cn/    http://www.int.ht0431.cn/    http://www.oqi.httx341.cn/    http://www.xhq.jfmjl45.cn/    http://www.o8g.jfoexx9.cn/    http://www.v2m.jlbyby120.cn/    http://www.kv6.jlxiehe.cn/    http://www.ki6.jzss412.cn/    http://www.3ti.lfbb172.cn/    http://www.i5j.nuxtf69.cn/    http://www.b7a.oiwrlk7.cn/    http://www.6ip.ovpiq76.cn/    http://www.yjv.piuye.cn/    http://www.6zm.pndd600.cn/    http://www.bhu.pwtkcj1.cn/    http://www.uym.qytag.cn/    http://www.hyo.rsbw019.cn/    http://www.y8h.shenbing120.cn/    http://www.21i.shenbingke120.cn/    http://www.8wx.shengbingke120.cn/    http://www.g4j.shenneike120.cn/    http://www.cgn.skdmc.cn/    http://www.15r.smzx120.cn/    http://www.vw0.swfq049.cn/    http://www.yzo.szbyy120.cn/    http://www.y7z.szqxe03.cn/    http://www.yja.thykd.cn/    http://www.z2f.tnaz800.cn/    http://www.7eq.tuphe.cn/    http://www.hpk.tyurk.cn/    http://www.lay.uyuhk.cn/    http://www.yd5.vmvq435.cn/    http://www.5c2.wdfgh.cn/    http://www.pyn.wiomh.cn/    http://www.yov.wjsk1199.cn/    http://www.qns.wjyy0431.cn/    http://www.ftc.wjyy1199.cn/    http://www.h70.woiti63.cn/    http://www.3d7.wulis.cn/    http://www.bfq.xbuh494.cn/    http://www.vhe.xhyy120.cn/    http://www.miq.ycestm1.cn/    http://www.w4v.ydy120.cn/    http://www.4sl.ygfk120.cn/    http://www.l98.ygrl120.cn/    http://www.5pa.ypjun54.cn/    http://www.7or.zafc120.cn/    http://www.egm.afygi.cn/    http://www.jw2.btexr.cn/    http://www.r9v.cznsu.cn/    http://www.xog.dmldf.cn/    http://www.xs4.jznzp.cn/    http://www.fev.pbcza.cn/    http://www.lov.udltv.cn/    http://www.6z5.urbxn.cn/    http://www.429.vjehn.cn/    http://www.2df.0431rl.cn/    http://www.h3u.0431wjyy.cn/    http://www.x6q.120girl.cn/    http://www.t5j.120shenbingke.cn/    http://www.rgi.120shenneike.cn/    http://www.jeg.120szbyy.cn/    http://www.v1k.120wjyy39.cn/    http://www.fi6.208fukew.cn/    http://www.hqr.521jk.cn/    http://www.23g.52fkw.cn/    http://www.ikf.********.cn/    http://www.ei2.********.cn/    http://www.q7b.********.cn/    http://www.rji.********.cn/    http://www.2f9.********.cn/    http://www.vwu.********.cn/    http://www.s2h.********.cn/    http://www.***-****1199.cn/    http://www.bnl.asqnf.cn/    http://www.isz.buyun365.cn/    http://www.1wq.bzhvcj4.cn/    http://www.qry.cc516.cn/    http://www.wym.ccby120.cn/    http://www.sn0.ccbyby.cn/    http://www.3t5.ccfk120.cn/    http://www.kz8.ccfkyy.cn/    http://www.1go.ccfkyy120.cn/    http://www.dv3.ccfuke.cn/    http://www.3ym.ccfuke120.cn/    http://www.6ud.cchmfk.cn/    http://www.vz6.ccmly120.cn/    http://www.mpy.ccrenliu.cn/    http://www.w5d.ccrl120.cn/    http://www.n4t.ccrlyy.cn/    http://www.97w.ccrsfk.cn/    http://www.534.ccsfuchan.cn/    http://www.j5w.ccshenbing120.cn/    http://www.0de.ccshenbing39.cn/    http://www.41b.ccszbyy120.cn/    http://www.kv8.ccwtrl.cn/    http://www.4jz.ccxhfk.cn/    http://www.50p.ccyc120.cn/    http://www.vb2.ccyg120.cn/    http://www.h4s.ccygfk.cn/    http://www.1vo.ccygfk120.cn/    http://www.k8d.ccygyy.cn/    http://www.jm9.ccygyy120.cn/    http://www.j57.dbbyby.cn/    http://www.isc.dslr120.cn/    http://www.hn5.eapaz36.cn/    http://www.3oq.fkylw.cn/    http://www.d9o.fkzx120.cn/    http://www.z6m.flxfd04.cn/    http://www.geq.gawga68.cn/    http://www.nc4.gmxlg45.cn/    http://www.vjn.gsofg48.cn/    http://www.zpj.gwy120.cn/    http://www.e9a.hmfk120.cn/    http://www.uza.ht0431.cn/    http://www.a4x.httx341.cn/    http://www.4bi.jfmjl45.cn/    http://www.ygw.jfoexx9.cn/    http://www.0qp.jlbyby120.cn/    http://www.a3n.jlxiehe.cn/    http://www.hsp.jzss412.cn/    http://www.k5b.lfbb172.cn/    http://www.9eq.nuxtf69.cn/    http://www.f43.oiwrlk7.cn/    http://www.bd6.ovpiq76.cn/    http://www.d3t.piuye.cn/    http://www.fw1.pndd600.cn/    http://www.7q8.pwtkcj1.cn/    http://www.pnt.qytag.cn/    http://www.7w8.rsbw019.cn/    http://www.d2m.shenbing120.cn/    http://www.2vx.shenbingke120.cn/    http://www.xjh.shengbingke120.cn/    http://www.fzb.shenneike120.cn/    http://www.gyv.skdmc.cn/    http://www.v92.smzx120.cn/    http://www.df3.swfq049.cn/    http://www.sep.szbyy120.cn/    http://www.16e.szqxe03.cn/    http://www.4t5.thykd.cn/    http://www.9l5.tnaz800.cn/    http://www.4if.tuphe.cn/    http://www.71u.tyurk.cn/    http://www.nl9.uyuhk.cn/    http://www.2j9.vmvq435.cn/    http://www.bp8.wdfgh.cn/    http://www.fb9.wiomh.cn/    http://www.31v.wjsk1199.cn/    http://www.yqe.wjyy0431.cn/    http://www.s0f.wjyy1199.cn/    http://www.1z6.woiti63.cn/    http://www.opk.wulis.cn/    http://www.uhv.xbuh494.cn/    http://www.pwk.xhyy120.cn/    http://www.hrt.ycestm1.cn/    http://www.7z3.ydy120.cn/    http://www.7k5.ygfk120.cn/    http://www.ezn.ygrl120.cn/    http://www.sdc.ypjun54.cn/    http://www.v78.zafc120.cn/    http://www.oxh.afygi.cn/    http://www.3i4.btexr.cn/    http://www.b9o.cznsu.cn/    http://www.8r2.dmldf.cn/    http://www.elr.jznzp.cn/    http://www.owv.pbcza.cn/    http://www.bhw.udltv.cn/    http://www.cp0.urbxn.cn/    http://www.9rd.vjehn.cn/    http://www.uw0.0431rl.cn/    http://www.4ux.0431wjyy.cn/    http://www.s3f.120girl.cn/    http://www.7wb.120shenbingke.cn/    http://www.c3b.120shenneike.cn/    http://www.yjr.120szbyy.cn/    http://www.4c3.120wjyy39.cn/    http://www.lm5.208fukew.cn/    http://www.lcm.521jk.cn/    http://www.bfj.52fkw.cn/    http://www.8va.********.cn/    http://www.kf5.********.cn/    http://www.n72.********.cn/    http://www.hov.********.cn/    http://www.d5g.********.cn/    http://www.xeb.********.cn/    http://www.v2e.********.cn/    http://www.ciy.********.cn/    http://www.ms4.asqnf.cn/    http://www.j62.buyun365.cn/    http://www.d83.bzhvcj4.cn/    http://www.13r.cc516.cn/    http://www.4zd.ccby120.cn/    http://www.gpb.ccbyby.cn/    http://www.xod.ccfk120.cn/    http://www.cvk.ccfkyy.cn/    http://www.jfb.ccfkyy120.cn/    http://www.kr1.ccfuke.cn/    http://www.7lt.ccfuke120.cn/    http://www.k7i.cchmfk.cn/    http://www.g65.ccmly120.cn/    http://www.lsp.ccrenliu.cn/    http://www.oxi.ccrl120.cn/    http://www.iuw.ccrlyy.cn/    http://www.7kc.ccrsfk.cn/    http://www.7h2.ccsfuchan.cn/    http://www.k3j.ccshenbing120.cn/    http://www.56p.ccshenbing39.cn/    http://www.ez5.ccszbyy120.cn/    http://www.1cg.ccwtrl.cn/    http://www.lwy.ccxhfk.cn/    http://www.ur5.ccyc120.cn/    http://www.kz7.ccyg120.cn/    http://www.9qh.ccygfk.cn/    http://www.4td.ccygfk120.cn/    http://www.yrs.ccygyy.cn/    http://www.5rb.ccygyy120.cn/    http://www.3i7.dbbyby.cn/    http://www.9d1.dslr120.cn/    http://www.w65.eapaz36.cn/    http://www.9fy.fkylw.cn/    http://www.xzj.fkzx120.cn/    http://www.blm.flxfd04.cn/    http://www.w5i.gawga68.cn/    http://www.bog.gmxlg45.cn/    http://www.p9w.gsofg48.cn/    http://www.gxj.gwy120.cn/    http://www.8su.hmfk120.cn/    http://www.sqz.ht0431.cn/    http://www.o76.httx341.cn/    http://www.4h0.jfmjl45.cn/    http://www.o4u.jfoexx9.cn/    http://www.zav.jlbyby120.cn/    http://www.yk0.jlxiehe.cn/    http://www.nyh.jzss412.cn/    http://www.p6b.lfbb172.cn/    http://www.yjt.nuxtf69.cn/    http://www.xhu.oiwrlk7.cn/    http://www.scj.ovpiq76.cn/    http://www.07r.piuye.cn/    http://www.3mc.pndd600.cn/    http://www.azv.pwtkcj1.cn/    http://www.mz9.qytag.cn/    http://www.lag.rsbw019.cn/    http://www.xko.shenbing120.cn/    http://www.1nr.shenbingke120.cn/    http://www.b02.shengbingke120.cn/    http://www.ws4.shenneike120.cn/    http://www.1hg.skdmc.cn/    http://www.kn1.smzx120.cn/    http://www.oax.swfq049.cn/    http://www.tyu.szbyy120.cn/    http://www.mpd.szqxe03.cn/    http://www.4dh.thykd.cn/    http://www.ehn.tnaz800.cn/    http://www.3ht.tuphe.cn/    http://www.l8m.tyurk.cn/    http://www.kgo.uyuhk.cn/    http://www.emx.vmvq435.cn/    http://www.b0y.wdfgh.cn/    http://www.z0b.wiomh.cn/    http://www.yn1.wjsk1199.cn/    http://www.zkg.wjyy0431.cn/    http://www.eiu.wjyy1199.cn/    http://www.2zi.woiti63.cn/    http://www.5oy.wulis.cn/    http://www.z46.xbuh494.cn/    http://www.98i.xhyy120.cn/    http://www.sj3.ycestm1.cn/    http://www.be6.ydy120.cn/    http://www.5f8.ygfk120.cn/    http://www.at8.ygrl120.cn/    http://www.7va.ypjun54.cn/    http://www.6aj.zafc120.cn/    http://www.lj9.afygi.cn/    http://www.r12.btexr.cn/    http://www.pyz.cznsu.cn/    http://www.z06.dmldf.cn/    http://www.xri.jznzp.cn/    http://www.dyu.pbcza.cn/    http://www.2wb.udltv.cn/    http://www.zl7.urbxn.cn/    http://www.no7.vjehn.cn/    http://www.hon.0431rl.cn/    http://www.ei5.0431wjyy.cn/    http://www.fms.120girl.cn/    http://www.qh3.120shenbingke.cn/    http://www.tuc.120shenneike.cn/    http://www.8tc.120szbyy.cn/    http://www.uyp.120wjyy39.cn/    http://www.04x.208fukew.cn/    http://www.dmk.521jk.cn/    http://www.vwm.52fkw.cn/    http://www.8hl.********.cn/    http://www.lin.********.cn/    http://www.04f.********.cn/    http://www.01r.********.cn/    http://www.o4y.********.cn/    http://www.n0x.********.cn/    http://www.63v.********.cn/    http://www.m39.********.cn/    http://www.e1c.asqnf.cn/    http://www.ec1.buyun365.cn/    http://www.now.bzhvcj4.cn/    http://www.jmi.cc516.cn/    http://www.gto.ccby120.cn/    http://www.75v.ccbyby.cn/    http://www.jlg.ccfk120.cn/    http://www.wfq.ccfkyy.cn/    http://www.39n.ccfkyy120.cn/    http://www.dtw.ccfuke.cn/    愿与食人野兽同流合污 可怜庇护于神殿之下的数百万南美幸存者绝对想不到 他们只是尊敬的神殿圣子口中之食。            “上次你做的过分了 不应该当面动手 至少不应该在没有确定弗兰德被杀死之前动手 现在我们还要面对弗兰德的报复 秘鲁和智利已经沦陷 丛林以每天三十公顷的面积消失 随着美国崩溃 越来越多的海族集中到南美 下个月丛林消失的速度也许会达到三百公顷 我们没有进化者 没有军队 甚至没有任何抵抗的能力 一旦南美沦陷 我们将无处藏身 你每天需要的十只羔羊也会断掉……。”|http://bbs.ent.163.com/bbs/bagua/605229403.html|2016-04-09
기타|2376397963|163_bbs|网易文化论坛-超级爆料|ZHO|2016-04-09 17:09:01|“那你有机会了 中国人准备突袭|大长老语气严肃起来 圣子并不在意 好看的眉毛轻挑 碧红的双眼闪动着玩味儿的光泽 扬起下巴说道：“那不是更好 我们到赤藻去藏身 每天享受高等海族的血肉不是更好？我的力量已经强大到无视高阶海族的地步 庇护数万人在赤藻生存没有问题 只要我和我的仆人们能像寄生虫那样吸食血族鲜血 就算地球毁灭了又有什么关系呢？上次击杀弗兰德的目的就是为了顶级进化者的血肉 我得到了就不算失败 等我能吞噬迪莉娅和厄俄斯 相信我会更加强大 像神一样强大……。”            大长老无奈的低下头 圣子生来与人类对立 这一点他很早就知道了 但他更知道想要得到永生和力量就必须和圣子合作 所以他出卖整个人类与圣子同流合污 但没想到圣子已经有了失去控制的迹象 让他心里也产生了微微的恐惧 南美洲并非一个进化者都没有 也许等圣子失去了最后的耐性 他这个曾经的第一使徒就会成为圣子的血食。http://www.a5e.woiti63.cn/    http://www.5kn.wulis.cn/    http://www.0iv.xbuh494.cn/    http://www.dws.xhyy120.cn/    http://www.t6m.ycestm1.cn/    http://www.xvo.ydy120.cn/    http://www.ydi.ygfk120.cn/    http://www.tzx.ygrl120.cn/    http://www.z1g.ypjun54.cn/    http://www.5oc.zafc120.cn/    http://www.u9o.afygi.cn/    http://www.6rh.btexr.cn/    http://www.mil.cznsu.cn/    http://www.vik.dmldf.cn/    http://www.7z6.jznzp.cn/    http://www.30x.pbcza.cn/    http://www.jet.udltv.cn/    http://www.sta.urbxn.cn/    http://www.et8.vjehn.cn/    http://www.28p.0431rl.cn/    http://www.p3w.0431wjyy.cn/    http://www.uoz.120girl.cn/    http://www.1sw.120shenbingke.cn/    http://www.4zf.120shenneike.cn/    http://www.uem.120szbyy.cn/    http://www.379.120wjyy39.cn/    http://www.yng.208fukew.cn/    http://www.u7j.521jk.cn/    http://www.1xc.52fkw.cn/    http://www.h2d.********.cn/    http://www.p5a.********.cn/    http://www.faw.********.cn/    http://www.0ma.********.cn/    http://www.2xz.********.cn/    http://www.cq4.********.cn/    http://www.bi0.********.cn/    http://www.bo3.********.cn/    http://www.fse.asqnf.cn/    http://www.cro.buyun365.cn/    http://www.2p4.bzhvcj4.cn/    http://www.4.00E+03.cc516.cn/    http://www.tfr.ccby120.cn/    http://www.gph.ccbyby.cn/    http://www.u2k.ccfk120.cn/    http://www.uhd.ccfkyy.cn/    http://www.nq7.ccfkyy120.cn/    http://www.iy3.ccfuke.cn/    http://www.qt3.ccfuke120.cn/    http://www.9wb.cchmfk.cn/    http://www.9c3.ccmly120.cn/    http://www.6zw.ccrenliu.cn/    http://www.17o.ccrl120.cn/    http://www.297.ccrlyy.cn/    http://www.az0.ccrsfk.cn/    http://www.md1.ccsfuchan.cn/    http://www.qlb.ccshenbing120.cn/    http://www.j0x.ccshenbing39.cn/    http://www.nh5.ccszbyy120.cn/    http://www.4of.ccwtrl.cn/    http://www.e82.ccxhfk.cn/    http://www.j8u.ccyc120.cn/    http://www.nbd.ccyg120.cn/    http://www.v7t.ccygfk.cn/    http://www.s9f.ccygfk120.cn/    http://www.e86.ccygyy.cn/    http://www.d6z.ccygyy120.cn/    http://www.i4u.dbbyby.cn/    http://www.ufe.dslr120.cn/    http://www.68j.eapaz36.cn/    http://www.01x.fkylw.cn/    http://www.6g3.fkzx120.cn/    http://www.kp5.flxfd04.cn/    http://www.si9.gawga68.cn/    http://www.xjb.gmxlg45.cn/    http://www.n8k.gsofg48.cn/    http://www.q8a.gwy120.cn/    http://www.47b.hmfk120.cn/    http://www.xwu.ht0431.cn/    http://www.ap8.httx341.cn/    http://www.hpk.jfmjl45.cn/    http://www.nlq.jfoexx9.cn/    http://www.m50.jlbyby120.cn/    http://www.ijz.jlxiehe.cn/    http://www.a8h.jzss412.cn/    http://www.ser.lfbb172.cn/    http://www.gpa.nuxtf69.cn/    http://www.g6e.oiwrlk7.cn/    http://www.2fm.ovpiq76.cn/    http://www.1jq.piuye.cn/    http://www.zd0.pndd600.cn/    http://www.y18.pwtkcj1.cn/    http://www.rh0.qytag.cn/    http://www.ftv.rsbw019.cn/    http://www.jap.shenbing120.cn/    http://www.q0p.shenbingke120.cn/    http://www.qhv.shengbingke120.cn/    http://www.59w.shenneike120.cn/    http://www.ukt.skdmc.cn/    http://www.jfo.smzx120.cn/    http://www.3wd.swfq049.cn/    http://www.mvb.szbyy120.cn/    http://www.lfi.szqxe03.cn/    http://www.9to.thykd.cn/    http://www.9x6.tnaz800.cn/    http://www.r7j.tuphe.cn/    http://www.d1l.tyurk.cn/    http://www.sy2.uyuhk.cn/    http://www.grz.vmvq435.cn/    http://www.my9.wdfgh.cn/    http://www.9ht.wiomh.cn/    http://www.cmg.wjsk1199.cn/    http://www.yus.wjyy0431.cn/    http://www.92y.wjyy1199.cn/    http://www.mht.woiti63.cn/    http://www.6zg.wulis.cn/    http://www.g10.xbuh494.cn/    http://www.cs6.xhyy120.cn/    http://www.ycs.ycestm1.cn/    http://www.9bz.ydy120.cn/    http://www.gfr.ygfk120.cn/    http://www.amc.ygrl120.cn/    http://www.fcq.ypjun54.cn/    http://www.key.zafc120.cn/    http://www.v0g.afygi.cn/    http://www.ruy.btexr.cn/    http://www.v0y.cznsu.cn/    http://www.tmf.dmldf.cn/    http://www.4ln.jznzp.cn/    http://www.rmc.pbcza.cn/    http://www.fji.udltv.cn/    http://www.98e.urbxn.cn/    http://www.8wa.vjehn.cn/    http://www.fkl.0431rl.cn/    http://www.e29.0431wjyy.cn/    http://www.4vj.120girl.cn/    http://www.heo.120shenbingke.cn/    http://www.m0l.120shenneike.cn/    http://www.dz2.120szbyy.cn/    http://www.et8.120wjyy39.cn/    http://www.foe.208fukew.cn/    http://www.i98.521jk.cn/    http://www.5bd.52fkw.cn/    http://www.2zd.********.cn/    http://www.iw2.********.cn/    http://www.v48.********.cn/    http://www.nd6.********.cn/    http://www.gjx.********.cn/    http://www.49s.********.cn/    http://www.jx7.********.cn/    http://www.sil.********.cn/    http://www.9ca.asqnf.cn/    http://www.60x.buyun365.cn/    http://www.obs.bzhvcj4.cn/    http://www.asb.cc516.cn/    http://www.1we.ccby120.cn/    http://www.5ci.ccbyby.cn/    http://www.3ij.ccfk120.cn/    http://www.78d.ccfkyy.cn/    http://www.a8s.ccfkyy120.cn/    http://www.tzp.ccfuke.cn/    http://www.wyb.ccfuke120.cn/    http://www.i4d.cchmfk.cn/    http://www.ezi.ccmly120.cn/    http://www.23l.ccrenliu.cn/    http://www.bne.ccrl120.cn/    http://www.kq8.ccrlyy.cn/    http://www.iac.ccrsfk.cn/    http://www.hv5.ccsfuchan.cn/    http://www.v0f.ccshenbing120.cn/    http://www.rz2.ccshenbing39.cn/    http://www.1rw.ccszbyy120.cn/    http://www.8jn.ccwtrl.cn/    http://www.hei.ccxhfk.cn/    http://www.ux9.ccyc120.cn/    http://www.hwe.ccyg120.cn/    http://www.ze3.ccygfk.cn/    http://www.cyo.ccygfk120.cn/    http://www.jl5.ccygyy.cn/    http://www.4qj.ccygyy120.cn/    http://www.3i1.dbbyby.cn/    http://www.u34.dslr120.cn/    http://www.28w.eapaz36.cn/    http://www.3lx.fkylw.cn/    http://www.du3.fkzx120.cn/    http://www.qif.flxfd04.cn/    http://www.ry1.gawga68.cn/    http://www.ul5.gmxlg45.cn/    http://www.nhv.gsofg48.cn/    http://www.f5x.gwy120.cn/    http://www.lue.hmfk120.cn/    http://www.int.ht0431.cn/    http://www.oqi.httx341.cn/    http://www.xhq.jfmjl45.cn/    http://www.o8g.jfoexx9.cn/    http://www.v2m.jlbyby120.cn/    http://www.kv6.jlxiehe.cn/    http://www.ki6.jzss412.cn/    http://www.3ti.lfbb172.cn/    http://www.i5j.nuxtf69.cn/    http://www.b7a.oiwrlk7.cn/    http://www.6ip.ovpiq76.cn/    http://www.yjv.piuye.cn/    http://www.6zm.pndd600.cn/    http://www.bhu.pwtkcj1.cn/    http://www.uym.qytag.cn/    http://www.hyo.rsbw019.cn/    http://www.y8h.shenbing120.cn/    http://www.21i.shenbingke120.cn/    http://www.8wx.shengbingke120.cn/    http://www.g4j.shenneike120.cn/    http://www.cgn.skdmc.cn/    http://www.15r.smzx120.cn/    http://www.vw0.swfq049.cn/    http://www.yzo.szbyy120.cn/    http://www.y7z.szqxe03.cn/    http://www.yja.thykd.cn/    http://www.z2f.tnaz800.cn/    http://www.7eq.tuphe.cn/    http://www.hpk.tyurk.cn/    http://www.lay.uyuhk.cn/    http://www.yd5.vmvq435.cn/    http://www.5c2.wdfgh.cn/    http://www.pyn.wiomh.cn/    http://www.yov.wjsk1199.cn/    http://www.qns.wjyy0431.cn/    http://www.ftc.wjyy1199.cn/    http://www.h70.woiti63.cn/    http://www.3d7.wulis.cn/    http://www.bfq.xbuh494.cn/    http://www.vhe.xhyy120.cn/    http://www.miq.ycestm1.cn/    http://www.w4v.ydy120.cn/    http://www.4sl.ygfk120.cn/    http://www.l98.ygrl120.cn/    http://www.5pa.ypjun54.cn/    http://www.7or.zafc120.cn/    http://www.egm.afygi.cn/    http://www.jw2.btexr.cn/    http://www.r9v.cznsu.cn/    http://www.xog.dmldf.cn/    http://www.xs4.jznzp.cn/    http://www.fev.pbcza.cn/    http://www.lov.udltv.cn/    http://www.6z5.urbxn.cn/    http://www.429.vjehn.cn/    http://www.2df.0431rl.cn/    http://www.h3u.0431wjyy.cn/    http://www.x6q.120girl.cn/    http://www.t5j.120shenbingke.cn/    http://www.rgi.120shenneike.cn/    http://www.jeg.120szbyy.cn/    http://www.v1k.120wjyy39.cn/    http://www.fi6.208fukew.cn/    http://www.hqr.521jk.cn/    http://www.23g.52fkw.cn/    http://www.ikf.********.cn/    http://www.ei2.********.cn/    http://www.q7b.********.cn/    http://www.rji.********.cn/    http://www.2f9.********.cn/    http://www.vwu.********.cn/    http://www.s2h.********.cn/    http://www.***-****1199.cn/    http://www.bnl.asqnf.cn/    http://www.isz.buyun365.cn/    http://www.1wq.bzhvcj4.cn/    http://www.qry.cc516.cn/    http://www.wym.ccby120.cn/    http://www.sn0.ccbyby.cn/    http://www.3t5.ccfk120.cn/    http://www.kz8.ccfkyy.cn/    http://www.1go.ccfkyy120.cn/    http://www.dv3.ccfuke.cn/    http://www.3ym.ccfuke120.cn/    http://www.6ud.cchmfk.cn/    http://www.vz6.ccmly120.cn/    http://www.mpy.ccrenliu.cn/    http://www.w5d.ccrl120.cn/    http://www.n4t.ccrlyy.cn/    http://www.97w.ccrsfk.cn/    http://www.534.ccsfuchan.cn/    http://www.j5w.ccshenbing120.cn/    http://www.0de.ccshenbing39.cn/    http://www.41b.ccszbyy120.cn/    http://www.kv8.ccwtrl.cn/    http://www.4jz.ccxhfk.cn/    http://www.50p.ccyc120.cn/    http://www.vb2.ccyg120.cn/    http://www.h4s.ccygfk.cn/    http://www.1vo.ccygfk120.cn/    http://www.k8d.ccygyy.cn/    http://www.jm9.ccygyy120.cn/    http://www.j57.dbbyby.cn/    http://www.isc.dslr120.cn/    http://www.hn5.eapaz36.cn/    http://www.3oq.fkylw.cn/    http://www.d9o.fkzx120.cn/    http://www.z6m.flxfd04.cn/    http://www.geq.gawga68.cn/    http://www.nc4.gmxlg45.cn/    http://www.vjn.gsofg48.cn/    http://www.zpj.gwy120.cn/    http://www.e9a.hmfk120.cn/    http://www.uza.ht0431.cn/    http://www.a4x.httx341.cn/    http://www.4bi.jfmjl45.cn/    http://www.ygw.jfoexx9.cn/    http://www.0qp.jlbyby120.cn/    http://www.a3n.jlxiehe.cn/    http://www.hsp.jzss412.cn/    http://www.k5b.lfbb172.cn/    http://www.9eq.nuxtf69.cn/    http://www.f43.oiwrlk7.cn/    http://www.bd6.ovpiq76.cn/    http://www.d3t.piuye.cn/    http://www.fw1.pndd600.cn/    http://www.7q8.pwtkcj1.cn/    http://www.pnt.qytag.cn/    http://www.7w8.rsbw019.cn/    http://www.d2m.shenbing120.cn/    http://www.2vx.shenbingke120.cn/    http://www.xjh.shengbingke120.cn/    http://www.fzb.shenneike120.cn/    http://www.gyv.skdmc.cn/    http://www.v92.smzx120.cn/    http://www.df3.swfq049.cn/    http://www.sep.szbyy120.cn/    http://www.16e.szqxe03.cn/    http://www.4t5.thykd.cn/    http://www.9l5.tnaz800.cn/    http://www.4if.tuphe.cn/    http://www.71u.tyurk.cn/    http://www.nl9.uyuhk.cn/    http://www.2j9.vmvq435.cn/    http://www.bp8.wdfgh.cn/    http://www.fb9.wiomh.cn/    http://www.31v.wjsk1199.cn/    http://www.yqe.wjyy0431.cn/    http://www.s0f.wjyy1199.cn/    http://www.1z6.woiti63.cn/    http://www.opk.wulis.cn/    http://www.uhv.xbuh494.cn/    http://www.pwk.xhyy120.cn/    http://www.hrt.ycestm1.cn/    http://www.7z3.ydy120.cn/    http://www.7k5.ygfk120.cn/    http://www.ezn.ygrl120.cn/    http://www.sdc.ypjun54.cn/    http://www.v78.zafc120.cn/    http://www.oxh.afygi.cn/    http://www.3i4.btexr.cn/    http://www.b9o.cznsu.cn/    http://www.8r2.dmldf.cn/    http://www.elr.jznzp.cn/    http://www.owv.pbcza.cn/    http://www.bhw.udltv.cn/    http://www.cp0.urbxn.cn/    http://www.9rd.vjehn.cn/    http://www.uw0.0431rl.cn/    http://www.4ux.0431wjyy.cn/    http://www.s3f.120girl.cn/    http://www.7wb.120shenbingke.cn/    http://www.c3b.120shenneike.cn/    http://www.yjr.120szbyy.cn/    http://www.4c3.120wjyy39.cn/    http://www.lm5.208fukew.cn/    http://www.lcm.521jk.cn/    http://www.bfj.52fkw.cn/    http://www.8va.********.cn/    http://www.kf5.********.cn/    http://www.n72.********.cn/    http://www.hov.********.cn/    http://www.d5g.********.cn/    http://www.xeb.********.cn/    http://www.v2e.********.cn/    http://www.ciy.********.cn/    http://www.ms4.asqnf.cn/    http://www.j62.buyun365.cn/    http://www.d83.bzhvcj4.cn/    http://www.13r.cc516.cn/    http://www.4zd.ccby120.cn/    http://www.gpb.ccbyby.cn/    http://www.xod.ccfk120.cn/    http://www.cvk.ccfkyy.cn/    http://www.jfb.ccfkyy120.cn/    http://www.kr1.ccfuke.cn/    http://www.7lt.ccfuke120.cn/    http://www.k7i.cchmfk.cn/    http://www.g65.ccmly120.cn/    http://www.lsp.ccrenliu.cn/    http://www.oxi.ccrl120.cn/    http://www.iuw.ccrlyy.cn/    http://www.7kc.ccrsfk.cn/    http://www.7h2.ccsfuchan.cn/    http://www.k3j.ccshenbing120.cn/    http://www.56p.ccshenbing39.cn/    http://www.ez5.ccszbyy120.cn/    http://www.1cg.ccwtrl.cn/    http://www.lwy.ccxhfk.cn/    http://www.ur5.ccyc120.cn/    http://www.kz7.ccyg120.cn/    http://www.9qh.ccygfk.cn/    http://www.4td.ccygfk120.cn/    http://www.yrs.ccygyy.cn/    http://www.5rb.ccygyy120.cn/    http://www.3i7.dbbyby.cn/    http://www.9d1.dslr120.cn/    http://www.w65.eapaz36.cn/    http://www.9fy.fkylw.cn/    http://www.xzj.fkzx120.cn/    http://www.blm.flxfd04.cn/    http://www.w5i.gawga68.cn/    http://www.bog.gmxlg45.cn/    http://www.p9w.gsofg48.cn/    http://www.gxj.gwy120.cn/    http://www.8su.hmfk120.cn/    http://www.sqz.ht0431.cn/    http://www.o76.httx341.cn/    http://www.4h0.jfmjl45.cn/    http://www.o4u.jfoexx9.cn/    http://www.zav.jlbyby120.cn/    http://www.yk0.jlxiehe.cn/    http://www.nyh.jzss412.cn/    http://www.p6b.lfbb172.cn/    http://www.yjt.nuxtf69.cn/    http://www.xhu.oiwrlk7.cn/    http://www.scj.ovpiq76.cn/    http://www.07r.piuye.cn/    http://www.3mc.pndd600.cn/    http://www.azv.pwtkcj1.cn/    http://www.mz9.qytag.cn/    http://www.lag.rsbw019.cn/    http://www.xko.shenbing120.cn/    http://www.1nr.shenbingke120.cn/    http://www.b02.shengbingke120.cn/    http://www.ws4.shenneike120.cn/    http://www.1hg.skdmc.cn/    http://www.kn1.smzx120.cn/    http://www.oax.swfq049.cn/    http://www.tyu.szbyy120.cn/    http://www.mpd.szqxe03.cn/    http://www.4dh.thykd.cn/    http://www.ehn.tnaz800.cn/    http://www.3ht.tuphe.cn/    http://www.l8m.tyurk.cn/    http://www.kgo.uyuhk.cn/    http://www.emx.vmvq435.cn/    http://www.b0y.wdfgh.cn/    http://www.z0b.wiomh.cn/    http://www.yn1.wjsk1199.cn/    http://www.zkg.wjyy0431.cn/    http://www.eiu.wjyy1199.cn/    http://www.2zi.woiti63.cn/    http://www.5oy.wulis.cn/    http://www.z46.xbuh494.cn/    http://www.98i.xhyy120.cn/    http://www.sj3.ycestm1.cn/    http://www.be6.ydy120.cn/    http://www.5f8.ygfk120.cn/    http://www.at8.ygrl120.cn/    http://www.7va.ypjun54.cn/    http://www.6aj.zafc120.cn/    http://www.lj9.afygi.cn/    http://www.r12.btexr.cn/    http://www.pyz.cznsu.cn/    http://www.z06.dmldf.cn/    http://www.xri.jznzp.cn/    http://www.dyu.pbcza.cn/    http://www.2wb.udltv.cn/    http://www.zl7.urbxn.cn/    http://www.no7.vjehn.cn/    http://www.hon.0431rl.cn/    http://www.ei5.0431wjyy.cn/    http://www.fms.120girl.cn/    http://www.qh3.120shenbingke.cn/    http://www.tuc.120shenneike.cn/    http://www.8tc.120szbyy.cn/    http://www.uyp.120wjyy39.cn/    http://www.04x.208fukew.cn/    http://www.dmk.521jk.cn/    http://www.vwm.52fkw.cn/    http://www.8hl.********.cn/    http://www.lin.********.cn/    http://www.04f.********.cn/    http://www.01r.********.cn/    http://www.o4y.********.cn/    http://www.n0x.********.cn/    http://www.63v.********.cn/    http://www.m39.********.cn/    http://www.e1c.asqnf.cn/    http://www.ec1.buyun365.cn/    http://www.now.bzhvcj4.cn/    http://www.jmi.cc516.cn/    http://www.gto.ccby120.cn/    http://www.75v.ccbyby.cn/    http://www.jlg.ccfk120.cn/    http://www.wfq.ccfkyy.cn/    http://www.39n.ccfkyy120.cn/    http://www.dtw.ccfuke.cn/    夏威夷海域 他们有能打破空中封锁的方法 迪莉娅和厄俄斯已经确定出动 中国人也有比他们不差的顶尖进化者出动……。”也许是因为害怕 也许是因为圣子已经超出了他的控制范围之外 大长老终于将这条消息说了出来。            “陷阱？”圣子用手指夹起餐刀在餐盘红白相间的肉块中翻动 那双敏感而纯净的眼睛却在偷偷扫视大元老。|http://bbs.ent.163.com/bbs/bagua/605229605.html|2016-04-09
其他媒体|2388686317|youku|生活|ZHO|2016-04-16 09:02:01|比亚迪S7遇小三前辈惊魂一幕||http://v.youku.com/v_show/id_XMTUzNjA3MTk3Mg==.html|2016-04-16
其他媒体|2389011980|zhidao_baidu|电脑/网络|ZHO|2016-04-16 13:51:01|海安那里有东风悦达起亚k3汽车车套买|汽车海安那里有东风悦达起亚k3汽车车套买|http://zhidao.baidu.com/question/875248707785204492.html?fr=qlquick&entry=qb_list_default|2016-04-16
其他媒体|2391070718|zhidao_baidu|电脑/网络 > 硬件 > 硬盘|ZHO|2016-04-17 21:39:01|起亚k3和广汽本田sus哪个好使用性更好|汽车起亚k3和广汽本田sus哪个好使用性更好|http://zhidao.baidu.com/question/714016742482089805.html?fr=qlquick&entry=qb_list_default|2016-04-17
其他媒体|2391073303|zhidao_baidu|烦恼|ZHO|2016-04-17 21:41:01|起亚k3和广汽本田sus哪个使用性更好|汽车起亚k3和广汽本田sus哪个使用性更好|http://zhidao.baidu.com/question/2269180814339904188.html?fr=qlquick&entry=qb_list_default|2016-04-17
기타|2415561013|Autohome review|혼다 어코드(雅阁)|ZHO|2016-04-30 17:26:02|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=107&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-04-30
기타|2415633648|Autohome review|혼다 어코드(雅阁)|ZHO|2016-04-30 18:22:03|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=108&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-04-30
기타|2415715277|Autohome review|혼다 어코드(雅阁)|ZHO|2016-04-30 19:24:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=109&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-04-30
기타|2415962653|Autohome review|혼다 어코드(雅阁)|ZHO|2016-04-30 22:37:04|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=110&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-04-30
기타|2418148448|Autohome review|혼다 어코드(雅阁)|ZHO|2016-05-02 10:19:02|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=115&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-02
기타|2418998456|Autohome review|혼다 어코드(雅阁)|ZHO|2016-05-02 19:02:02|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=116&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-02
기타|2419436432|Autohome review|혼다 어코드(雅阁)|ZHO|2016-05-02 23:45:02|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=117&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-02
기타|2464972009|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 00:21:07|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=173&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2464975488|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-27 00:24:05|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=142&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-27
其他媒体|2464990354|bitauto|易车 > 问答 > 问题分类|ZHO|2016-05-27 00:35:02|雷凌包真皮好吗？4s报价2500是真皮吗？我的是精英版 原车|雷凌包真皮好吗？4s报价2500是真皮吗？我的是精英版 原车     提问者：伤逝k38y6o  分类：  丰田  雷凌  买车  车型  浏览[8] 来自：易车手机客户端  2016-05-26 23:24  举报   雷凌包真皮好吗？4s报价2500是真皮吗？我的是精英版 原车配的是织物|http://ask.bitauto.com/detail/6595850/?leads_source=p029001|2016-05-27
기타|2465021699|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-27 00:54:01|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=141&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-27
기타|2465023628|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 00:55:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=154&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2465023759|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 00:55:01|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=110&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-27
기타|2465034045|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-27 01:02:02|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=201&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-27
기타|2465076080|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-27 01:34:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=101&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2465087154|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 01:42:01|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=105&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-27
기타|2465087323|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 01:42:01|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=46&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-27
기타|2465100748|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 01:54:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=155&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2465100841|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 01:54:01|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=111&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-27
기타|2465109842|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-27 02:02:01|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=203&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-27
기타|2465118773|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 02:09:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=174&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2465144248|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-27 02:35:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=102&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2465154783|Autohome_review|랑동(朗动)|ZHO|2016-05-27 02:45:01|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=172&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-27
기타|2465172785|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 03:06:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=176&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2465198196|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 03:36:01|2016年04月23日 发表了口碑|来自：手机汽车之家  2016年04月23日 发表了口碑  口碑    《外形流线、内饰满意 油耗经济 钣金太薄 基本满意》             【最满意的一点】最满意的就是整体车的线条和内饰 动力方面家用足够了、油耗方面觉得比较省油 目前油耗7.2._7.9。磨合完了可能还能降低 方向很轻 指向性还是不错的 空间方面也比较满意 后排中间是平的 日韩好象都这样 后排中间靠背可以放下来当杯架和扶手 和后备箱是通的 这个还是比较方便。有esp加前后气囊 再加开车时候遵守交通规则 多少也能弥补钣金薄的缺点 总体还是比较满意的【最不满意的一点】钣金太薄 后备箱盖子薄的就像饼干桶 中控有点塑料感 大灯角度调节形同虚设 大灯的亮度不够 有车友用蜡烛灯来比喻 其他还没发现【空间】【动力】电脑分配延迟大概一秒【操控】方向轻 指向性还是不错的【油耗】75的油耗不算费油【舒适性】启动和30码以内真心静音 80码以上开始胎噪有点大【外观】这个外观是满意的【内饰】基本满意【性价比】家用车中性价比还算不错 外观 油耗 空间都能4分以上。钣金、钣金 钣金    你门懂得。每个人心中自己的车是不一样的 我也就是在这里谈谈自己的感受。目前才500公里、首保后再和大家分享下感受【为什么最终选择这款车？】其实当时买车没考虑这款 朗行和卡罗拉是我的首选、路过起亚店 一见钟情型吧、就选中了16款k3、我个人消费能力之内随意性比较大、销售灰常的热情 我也觉得16款外形 内饰 油耗 内饰也是我预算范围内的 就小卡一刷【其他描述】改装中 内饰装修 车顶膜 大灯|http://k.autohome.com.cn/spec/19724/view_1084435_1.html?st=186&piap=0 2886 0 0 2 0 0 0 0 0 1#20160423|2016-05-27
기타|2465198236|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 03:36:01|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=168&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-05-27
기타|2465198464|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 03:36:01|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=84&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-05-27
기타|2465198493|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 03:36:01|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。【最不满意的一点】买的自动挡的 动力比较弱 超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 隔音也不咋地 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 本来就打算定福睿斯了 51和姐夫一起去车展看福睿斯的 姐夫说福睿斯不咋地 屁股太丑 16款的k3还不错 然后我就考虑了一下 就定了k3 因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的。|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=66&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-05-27
기타|2465198496|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 03:36:01|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=63&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-05-27
기타|2465198682|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 03:36:01|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=107&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-27
기타|2465198789|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 03:36:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=48&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-27
기타|2465241647|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 04:39:03|2016年04月23日 发表了口碑|来自：手机汽车之家  2016年04月23日 发表了口碑  口碑    《外形流线、内饰满意 油耗经济 钣金太薄 基本满意》             【最满意的一点】最满意的就是整体车的线条和内饰 动力方面家用足够了、油耗方面觉得比较省油 目前油耗7.2._7.9。磨合完了可能还能降低 方向很轻 指向性还是不错的 空间方面也比较满意 后排中间是平的 日韩好象都这样 后排中间靠背可以放下来当杯架和扶手 和后备箱是通的 这个还是比较方便。有esp加前后气囊 再加开车时候遵守交通规则 多少也能弥补钣金薄的缺点 总体还是比较满意的【最不满意的一点】钣金太薄 后备箱盖子薄的就像饼干桶 中控有点塑料感 大灯角度调节形同虚设 大灯的亮度不够 有车友用蜡烛灯来比喻 其他还没发现【空间】【动力】电脑分配延迟大概一秒【操控】方向轻 指向性还是不错的【油耗】75的油耗不算费油【舒适性】启动和30码以内真心静音 80码以上开始胎噪有点大【外观】这个外观是满意的【内饰】基本满意【性价比】家用车中性价比还算不错 外观 油耗 空间都能4分以上。钣金、钣金 钣金    你门懂得。每个人心中自己的车是不一样的 我也就是在这里谈谈自己的感受。目前才500公里、首保后再和大家分享下感受【为什么最终选择这款车？】其实当时买车没考虑这款 朗行和卡罗拉是我的首选、路过起亚店 一见钟情型吧、就选中了16款k3、我个人消费能力之内随意性比较大、销售灰常的热情 我也觉得16款外形 内饰 油耗 内饰也是我预算范围内的 就小卡一刷【其他描述】改装中 内饰装修 车顶膜 大灯|http://k.autohome.com.cn/spec/19724/view_1084435_1.html?st=187&piap=0 2886 0 0 2 0 0 0 0 0 1#20160423|2016-05-27
기타|2465241711|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 04:39:03|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=169&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-05-27
기타|2465241893|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 04:39:03|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=85&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-05-27
기타|2465241933|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 04:39:03|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。【最不满意的一点】买的自动挡的 动力比较弱 超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 隔音也不咋地 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 本来就打算定福睿斯了 51和姐夫一起去车展看福睿斯的 姐夫说福睿斯不咋地 屁股太丑 16款的k3还不错 然后我就考虑了一下 就定了k3 因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的。|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=67&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-05-27
기타|2465241938|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 04:39:03|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=64&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-05-27
기타|2465243029|Autohome_review|랑동(朗动)|ZHO|2016-05-27 04:41:02|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=173&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-27
기타|2465353514|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 07:25:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=177&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2465353600|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 07:25:01|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=108&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-27
기타|2465353862|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 07:25:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=49&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-27
기타|2465492444|Autohome_review|랑동(朗动)|ZHO|2016-05-27 09:35:02|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=174&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-27
기타|2465577847|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-27 10:30:01|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=204&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-27
기타|2465584861|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-27 10:35:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=103&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2465690744|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 11:33:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=156&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2465690887|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 11:33:01|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=112&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-27
기타|2465713012|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-27 11:45:01|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=206&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-27
其他媒体|2465731370|bitauto|易车 > 问答 > 问题分类|ZHO|2016-05-27 11:55:03|东风悦达起亚k3 450公里多少油钱|东风悦达起亚k3 450公里多少油钱     提问者：易车网友 分类：  东风  二手车  评估  浏览[3]  2016-05-27 10:49  举报   东风悦达起亚k3 450公里多少油钱|http://ask.bitauto.com/detail/6596783/?leads_source=p029001|2016-05-27
기타|2465778985|Autohome_review|랑동(朗动)|ZHO|2016-05-27 12:22:02|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=175&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-27
기타|2465812604|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-27 12:44:02|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=208&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-27
기타|2465867369|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-27 13:20:17|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=105&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2465875676|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 13:25:16|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=159&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2465875733|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 13:25:16|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=115&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-27
기타|2465902633|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-27 13:43:01|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=209&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-27
기타|2465910629|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 13:48:01|2016年04月23日 发表了口碑|来自：手机汽车之家  2016年04月23日 发表了口碑  口碑    《外形流线、内饰满意 油耗经济 钣金太薄 基本满意》             【最满意的一点】最满意的就是整体车的线条和内饰 动力方面家用足够了、油耗方面觉得比较省油 目前油耗7.2._7.9。磨合完了可能还能降低 方向很轻 指向性还是不错的 空间方面也比较满意 后排中间是平的 日韩好象都这样 后排中间靠背可以放下来当杯架和扶手 和后备箱是通的 这个还是比较方便。有esp加前后气囊 再加开车时候遵守交通规则 多少也能弥补钣金薄的缺点 总体还是比较满意的【最不满意的一点】钣金太薄 后备箱盖子薄的就像饼干桶 中控有点塑料感 大灯角度调节形同虚设 大灯的亮度不够 有车友用蜡烛灯来比喻 其他还没发现【空间】【动力】电脑分配延迟大概一秒【操控】方向轻 指向性还是不错的【油耗】75的油耗不算费油【舒适性】启动和30码以内真心静音 80码以上开始胎噪有点大【外观】这个外观是满意的【内饰】基本满意【性价比】家用车中性价比还算不错 外观 油耗 空间都能4分以上。钣金、钣金 钣金    你门懂得。每个人心中自己的车是不一样的 我也就是在这里谈谈自己的感受。目前才500公里、首保后再和大家分享下感受【为什么最终选择这款车？】其实当时买车没考虑这款 朗行和卡罗拉是我的首选、路过起亚店 一见钟情型吧、就选中了16款k3、我个人消费能力之内随意性比较大、销售灰常的热情 我也觉得16款外形 内饰 油耗 内饰也是我预算范围内的 就小卡一刷【其他描述】改装中 内饰装修 车顶膜 大灯|http://k.autohome.com.cn/spec/19724/view_1084435_1.html?st=188&piap=0 2886 0 0 2 0 0 0 0 0 1#20160423|2016-05-27
기타|2465910688|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 13:48:01|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=170&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-05-27
기타|2465910886|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 13:48:01|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=86&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-05-27
기타|2465910914|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 13:48:01|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。【最不满意的一点】买的自动挡的 动力比较弱 超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 隔音也不咋地 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 本来就打算定福睿斯了 51和姐夫一起去车展看福睿斯的 姐夫说福睿斯不咋地 屁股太丑 16款的k3还不错 然后我就考虑了一下 就定了k3 因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的。|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=68&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-05-27
기타|2465910918|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 13:48:01|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=65&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-05-27
기타|2465917252|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-27 13:52:05|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=106&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2466005476|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 14:47:30|2016年04月23日 发表了口碑|来自：手机汽车之家  2016年04月23日 发表了口碑  口碑    《外形流线、内饰满意 油耗经济 钣金太薄 基本满意》             【最满意的一点】最满意的就是整体车的线条和内饰 动力方面家用足够了、油耗方面觉得比较省油 目前油耗7.2._7.9。磨合完了可能还能降低 方向很轻 指向性还是不错的 空间方面也比较满意 后排中间是平的 日韩好象都这样 后排中间靠背可以放下来当杯架和扶手 和后备箱是通的 这个还是比较方便。有esp加前后气囊 再加开车时候遵守交通规则 多少也能弥补钣金薄的缺点 总体还是比较满意的【最不满意的一点】钣金太薄 后备箱盖子薄的就像饼干桶 中控有点塑料感 大灯角度调节形同虚设 大灯的亮度不够 有车友用蜡烛灯来比喻 其他还没发现【空间】【动力】电脑分配延迟大概一秒【操控】方向轻 指向性还是不错的【油耗】75的油耗不算费油【舒适性】启动和30码以内真心静音 80码以上开始胎噪有点大【外观】这个外观是满意的【内饰】基本满意【性价比】家用车中性价比还算不错 外观 油耗 空间都能4分以上。钣金、钣金 钣金    你门懂得。每个人心中自己的车是不一样的 我也就是在这里谈谈自己的感受。目前才500公里、首保后再和大家分享下感受【为什么最终选择这款车？】其实当时买车没考虑这款 朗行和卡罗拉是我的首选、路过起亚店 一见钟情型吧、就选中了16款k3、我个人消费能力之内随意性比较大、销售灰常的热情 我也觉得16款外形 内饰 油耗 内饰也是我预算范围内的 就小卡一刷【其他描述】改装中 内饰装修 车顶膜 大灯|http://k.autohome.com.cn/spec/19724/view_1084435_1.html?st=189&piap=0 2886 0 0 2 0 0 0 0 0 1#20160423|2016-05-27
기타|2466005502|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 14:47:30|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=171&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-05-27
기타|2466006148|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 14:47:30|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=87&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-05-27
기타|2466006177|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 14:47:31|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。【最不满意的一点】买的自动挡的 动力比较弱 超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 隔音也不咋地 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 本来就打算定福睿斯了 51和姐夫一起去车展看福睿斯的 姐夫说福睿斯不咋地 屁股太丑 16款的k3还不错 然后我就考虑了一下 就定了k3 因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的。|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=69&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-05-27
기타|2466006180|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 14:47:31|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=66&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-05-27
기타|2466036201|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 15:07:22|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=179&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2466036287|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 15:07:22|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=110&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-27
기타|2466036357|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 15:07:22|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=51&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-27
기타|2466065798|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 15:28:29|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=162&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2466067507|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 15:28:38|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=118&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-27
기타|2466103841|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 15:46:10|2016年04月23日 发表了口碑|来自：手机汽车之家  2016年04月23日 发表了口碑  口碑    《外形流线、内饰满意 油耗经济 钣金太薄 基本满意》             【最满意的一点】最满意的就是整体车的线条和内饰 动力方面家用足够了、油耗方面觉得比较省油 目前油耗7.2._7.9。磨合完了可能还能降低 方向很轻 指向性还是不错的 空间方面也比较满意 后排中间是平的 日韩好象都这样 后排中间靠背可以放下来当杯架和扶手 和后备箱是通的 这个还是比较方便。有esp加前后气囊 再加开车时候遵守交通规则 多少也能弥补钣金薄的缺点 总体还是比较满意的【最不满意的一点】钣金太薄 后备箱盖子薄的就像饼干桶 中控有点塑料感 大灯角度调节形同虚设 大灯的亮度不够 有车友用蜡烛灯来比喻 其他还没发现【空间】【动力】电脑分配延迟大概一秒【操控】方向轻 指向性还是不错的【油耗】75的油耗不算费油【舒适性】启动和30码以内真心静音 80码以上开始胎噪有点大【外观】这个外观是满意的【内饰】基本满意【性价比】家用车中性价比还算不错 外观 油耗 空间都能4分以上。钣金、钣金 钣金    你门懂得。每个人心中自己的车是不一样的 我也就是在这里谈谈自己的感受。目前才500公里、首保后再和大家分享下感受【为什么最终选择这款车？】其实当时买车没考虑这款 朗行和卡罗拉是我的首选、路过起亚店 一见钟情型吧、就选中了16款k3、我个人消费能力之内随意性比较大、销售灰常的热情 我也觉得16款外形 内饰 油耗 内饰也是我预算范围内的 就小卡一刷【其他描述】改装中 内饰装修 车顶膜 大灯|http://k.autohome.com.cn/spec/19724/view_1084435_1.html?st=192&piap=0 2886 0 0 2 0 0 0 0 0 1#20160423|2016-05-27
기타|2466104051|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 15:46:10|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=174&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-05-27
기타|2466104583|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 15:46:11|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=90&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-05-27
기타|2466104658|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 15:46:11|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。【最不满意的一点】买的自动挡的 动力比较弱 超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 隔音也不咋地 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 本来就打算定福睿斯了 51和姐夫一起去车展看福睿斯的 姐夫说福睿斯不咋地 屁股太丑 16款的k3还不错 然后我就考虑了一下 就定了k3 因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的。|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=72&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-05-27
기타|2466104676|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 15:46:11|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=69&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-05-27
기타|2466124969|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 15:59:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=163&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2466125064|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 15:59:01|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=119&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-27
기타|2466190209|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-27 16:44:09|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=143&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-27
기타|2466191654|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-27 16:44:10|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=210&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-27
기타|2466205857|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 16:48:07|2016年04月23日 发表了口碑|来自：手机汽车之家  2016年04月23日 发表了口碑  口碑    《外形流线、内饰满意 油耗经济 钣金太薄 基本满意》             【最满意的一点】最满意的就是整体车的线条和内饰 动力方面家用足够了、油耗方面觉得比较省油 目前油耗7.2._7.9。磨合完了可能还能降低 方向很轻 指向性还是不错的 空间方面也比较满意 后排中间是平的 日韩好象都这样 后排中间靠背可以放下来当杯架和扶手 和后备箱是通的 这个还是比较方便。有esp加前后气囊 再加开车时候遵守交通规则 多少也能弥补钣金薄的缺点 总体还是比较满意的【最不满意的一点】钣金太薄 后备箱盖子薄的就像饼干桶 中控有点塑料感 大灯角度调节形同虚设 大灯的亮度不够 有车友用蜡烛灯来比喻 其他还没发现【空间】【动力】电脑分配延迟大概一秒【操控】方向轻 指向性还是不错的【油耗】75的油耗不算费油【舒适性】启动和30码以内真心静音 80码以上开始胎噪有点大【外观】这个外观是满意的【内饰】基本满意【性价比】家用车中性价比还算不错 外观 油耗 空间都能4分以上。钣金、钣金 钣金    你门懂得。每个人心中自己的车是不一样的 我也就是在这里谈谈自己的感受。目前才500公里、首保后再和大家分享下感受【为什么最终选择这款车？】其实当时买车没考虑这款 朗行和卡罗拉是我的首选、路过起亚店 一见钟情型吧、就选中了16款k3、我个人消费能力之内随意性比较大、销售灰常的热情 我也觉得16款外形 内饰 油耗 内饰也是我预算范围内的 就小卡一刷【其他描述】改装中 内饰装修 车顶膜 大灯|http://k.autohome.com.cn/spec/19724/view_1084435_1.html?st=193&piap=0 2886 0 0 2 0 0 0 0 0 1#20160423|2016-05-27
기타|2466205916|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 16:48:07|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=175&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-05-27
기타|2466207806|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 16:49:02|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=91&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-05-27
기타|2466207835|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 16:49:02|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。【最不满意的一点】买的自动挡的 动力比较弱 超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 隔音也不咋地 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 本来就打算定福睿斯了 51和姐夫一起去车展看福睿斯的 姐夫说福睿斯不咋地 屁股太丑 16款的k3还不错 然后我就考虑了一下 就定了k3 因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的。|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=73&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-05-27
기타|2466207839|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 16:49:02|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=70&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-05-27
기타|2466229585|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-27 16:57:03|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=107&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2466235972|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 17:01:01|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=120&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-27
기타|2466238801|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 17:02:01|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=111&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-27
기타|2466239208|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 17:02:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=52&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-27
기타|2466261939|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-27 17:16:03|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=145&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-27
기타|2466266395|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-27 17:19:12|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=212&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-27
기타|2466298181|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 17:35:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=181&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2466299495|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 17:36:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=164&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2466327083|Autohome_review|랑동(朗动)|ZHO|2016-05-27 17:51:01|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=176&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-27
기타|2466330302|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-27 17:53:02|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=213&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-27
기타|2466351299|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 18:04:01|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=112&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-27
기타|2466351398|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 18:04:01|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=53&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-27
기타|2466364953|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 18:12:09|2016年04月23日 发表了口碑|来自：手机汽车之家  2016年04月23日 发表了口碑  口碑    《外形流线、内饰满意 油耗经济 钣金太薄 基本满意》             【最满意的一点】最满意的就是整体车的线条和内饰 动力方面家用足够了、油耗方面觉得比较省油 目前油耗7.2._7.9。磨合完了可能还能降低 方向很轻 指向性还是不错的 空间方面也比较满意 后排中间是平的 日韩好象都这样 后排中间靠背可以放下来当杯架和扶手 和后备箱是通的 这个还是比较方便。有esp加前后气囊 再加开车时候遵守交通规则 多少也能弥补钣金薄的缺点 总体还是比较满意的【最不满意的一点】钣金太薄 后备箱盖子薄的就像饼干桶 中控有点塑料感 大灯角度调节形同虚设 大灯的亮度不够 有车友用蜡烛灯来比喻 其他还没发现【空间】【动力】电脑分配延迟大概一秒【操控】方向轻 指向性还是不错的【油耗】75的油耗不算费油【舒适性】启动和30码以内真心静音 80码以上开始胎噪有点大【外观】这个外观是满意的【内饰】基本满意【性价比】家用车中性价比还算不错 外观 油耗 空间都能4分以上。钣金、钣金 钣金    你门懂得。每个人心中自己的车是不一样的 我也就是在这里谈谈自己的感受。目前才500公里、首保后再和大家分享下感受【为什么最终选择这款车？】其实当时买车没考虑这款 朗行和卡罗拉是我的首选、路过起亚店 一见钟情型吧、就选中了16款k3、我个人消费能力之内随意性比较大、销售灰常的热情 我也觉得16款外形 内饰 油耗 内饰也是我预算范围内的 就小卡一刷【其他描述】改装中 内饰装修 车顶膜 大灯|http://k.autohome.com.cn/spec/19724/view_1084435_1.html?st=194&piap=0 2886 0 0 2 0 0 0 0 0 1#20160423|2016-05-27
기타|2466365000|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 18:12:09|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=176&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-05-27
기타|2466365188|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 18:12:09|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=92&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-05-27
기타|2466365236|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 18:12:09|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。【最不满意的一点】买的自动挡的 动力比较弱 超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 隔音也不咋地 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 本来就打算定福睿斯了 51和姐夫一起去车展看福睿斯的 姐夫说福睿斯不咋地 屁股太丑 16款的k3还不错 然后我就考虑了一下 就定了k3 因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的。|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=74&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-05-27
기타|2466365243|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 18:12:09|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=71&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-05-27
기타|2466390774|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-27 18:28:04|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=214&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-27
기타|2466411779|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 18:38:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=183&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2466412006|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 18:38:02|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=113&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-27
기타|2466412085|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 18:38:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=54&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-27
기타|2466428255|Autohome_review|랑동(朗动)|ZHO|2016-05-27 18:47:49|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=177&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-27
기타|2466461995|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 19:06:01|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=55&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-27
기타|2466471331|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-27 19:12:04|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=146&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-27
기타|2466491873|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-27 19:24:01|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=216&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-27
기타|2466507034|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 19:34:01|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=114&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-27
기타|2466553244|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 20:02:01|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=56&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-27
기타|2466560719|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 20:07:22|2016年04月23日 发表了口碑|来自：手机汽车之家  2016年04月23日 发表了口碑  口碑    《外形流线、内饰满意 油耗经济 钣金太薄 基本满意》             【最满意的一点】最满意的就是整体车的线条和内饰 动力方面家用足够了、油耗方面觉得比较省油 目前油耗7.2._7.9。磨合完了可能还能降低 方向很轻 指向性还是不错的 空间方面也比较满意 后排中间是平的 日韩好象都这样 后排中间靠背可以放下来当杯架和扶手 和后备箱是通的 这个还是比较方便。有esp加前后气囊 再加开车时候遵守交通规则 多少也能弥补钣金薄的缺点 总体还是比较满意的【最不满意的一点】钣金太薄 后备箱盖子薄的就像饼干桶 中控有点塑料感 大灯角度调节形同虚设 大灯的亮度不够 有车友用蜡烛灯来比喻 其他还没发现【空间】【动力】电脑分配延迟大概一秒【操控】方向轻 指向性还是不错的【油耗】75的油耗不算费油【舒适性】启动和30码以内真心静音 80码以上开始胎噪有点大【外观】这个外观是满意的【内饰】基本满意【性价比】家用车中性价比还算不错 外观 油耗 空间都能4分以上。钣金、钣金 钣金    你门懂得。每个人心中自己的车是不一样的 我也就是在这里谈谈自己的感受。目前才500公里、首保后再和大家分享下感受【为什么最终选择这款车？】其实当时买车没考虑这款 朗行和卡罗拉是我的首选、路过起亚店 一见钟情型吧、就选中了16款k3、我个人消费能力之内随意性比较大、销售灰常的热情 我也觉得16款外形 内饰 油耗 内饰也是我预算范围内的 就小卡一刷【其他描述】改装中 内饰装修 车顶膜 大灯|http://k.autohome.com.cn/spec/19724/view_1084435_1.html?st=195&piap=0 2886 0 0 2 0 0 0 0 0 1#20160423|2016-05-27
기타|2466560776|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 20:07:22|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=177&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-05-27
기타|2466560917|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 20:07:22|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=93&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-05-27
기타|2466560989|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 20:07:22|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。【最不满意的一点】买的自动挡的 动力比较弱 超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 隔音也不咋地 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 本来就打算定福睿斯了 51和姐夫一起去车展看福睿斯的 姐夫说福睿斯不咋地 屁股太丑 16款的k3还不错 然后我就考虑了一下 就定了k3 因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的。|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=75&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-05-27
기타|2466561001|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 20:07:22|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=72&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-05-27
기타|2466582225|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-27 20:20:03|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=217&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-27
기타|2466600781|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 20:32:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=184&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2466600929|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 20:32:02|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=115&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-27
기타|2466612592|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 20:39:02|2016年04月23日 发表了口碑|来自：手机汽车之家  2016年04月23日 发表了口碑  口碑    《外形流线、内饰满意 油耗经济 钣金太薄 基本满意》             【最满意的一点】最满意的就是整体车的线条和内饰 动力方面家用足够了、油耗方面觉得比较省油 目前油耗7.2._7.9。磨合完了可能还能降低 方向很轻 指向性还是不错的 空间方面也比较满意 后排中间是平的 日韩好象都这样 后排中间靠背可以放下来当杯架和扶手 和后备箱是通的 这个还是比较方便。有esp加前后气囊 再加开车时候遵守交通规则 多少也能弥补钣金薄的缺点 总体还是比较满意的【最不满意的一点】钣金太薄 后备箱盖子薄的就像饼干桶 中控有点塑料感 大灯角度调节形同虚设 大灯的亮度不够 有车友用蜡烛灯来比喻 其他还没发现【空间】【动力】电脑分配延迟大概一秒【操控】方向轻 指向性还是不错的【油耗】75的油耗不算费油【舒适性】启动和30码以内真心静音 80码以上开始胎噪有点大【外观】这个外观是满意的【内饰】基本满意【性价比】家用车中性价比还算不错 外观 油耗 空间都能4分以上。钣金、钣金 钣金    你门懂得。每个人心中自己的车是不一样的 我也就是在这里谈谈自己的感受。目前才500公里、首保后再和大家分享下感受【为什么最终选择这款车？】其实当时买车没考虑这款 朗行和卡罗拉是我的首选、路过起亚店 一见钟情型吧、就选中了16款k3、我个人消费能力之内随意性比较大、销售灰常的热情 我也觉得16款外形 内饰 油耗 内饰也是我预算范围内的 就小卡一刷【其他描述】改装中 内饰装修 车顶膜 大灯|http://k.autohome.com.cn/spec/19724/view_1084435_1.html?st=196&piap=0 2886 0 0 2 0 0 0 0 0 1#20160423|2016-05-27
기타|2466621671|Autohome_review|랑동(朗动)|ZHO|2016-05-27 20:44:03|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=178&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-27
기타|2466629702|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-27 20:51:01|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=219&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-27
기타|2466641231|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 20:58:03|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=165&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2466641370|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 20:58:03|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=121&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-27
기타|2466656655|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 21:07:25|2016年04月26日 发表了口碑|来自：手机汽车之家  2016年04月26日 发表了口碑  口碑   《这个价位的车性价比算高的了》   【最满意的一点】外观【最不满意的一点】低配差太多东西了 没有esp【空间】空间挺大 就是后排不能放倒有些遗憾【动力】起步很弱【操控】转向还好 就是路感很强【油耗】刚跑几天油耗就在八个多油了 挺好【舒适性】低配 你懂的【外观】喜欢这个设计【内饰】这个价位 内饰算好的了【性价比】如果有esp就给满分【为什么最终选择这款车？】实话实说选择这个车我自己都觉得很意外 之前家里人一直推荐卡罗拉但是本着些许爱国情节和极度不喜的内饰最终pass掉了 后来关注吉利博越上市后试驾了一次 感觉真是个好车 不管外观还是内饰都挺喜欢 要是吉利有免息金融贷款肯定就买了 可惜没有加上是新车没有接受市场的检验还是决定不当小白鼠了！九号看了苏州广电搞的车展没什么惊喜 回来在汽车之家搜了搜十万左右的车 偶然发现起亚k3优惠巨大 后来就买了它！【其他描述】|http://k.autohome.com.cn/spec/25737/view_1089742_1.html?st=178&piap=0 2886 0 0 2 0 0 0 0 0 1#20160426|2016-05-27
기타|2466656764|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 21:07:26|2016年05月10日 发表了口碑|来自：手机汽车之家  2016年05月10日 发表了口碑  口碑    《家用代步完全够用！酷酷的！》           【最满意的一点】外观拉风 酷酷的日间行车灯！油耗控制的非常好 省油！【最不满意的一点】起步时动力稍弱 真皮座椅 还有中控大屏还要选装！！【空间】后排空间稍小 前排还算够用【动力】起步就不谈了 除非给大油！跑起来就好多了 超车无压力！【操控】转向精准 只是过稍微颠簸路面的时候 车里不是很舒服 感觉不是那么稳！【油耗】油耗很满意 综合油耗7个！自动挡这个油耗真的是够省油的了！【舒适性】不是真皮座椅 套上了坐垫 感觉包裹性没有了！五一出了趟远门感觉不累！空调是真的很给力 很爽 非常舒服！只是后排没有空调口【外观】外观不说了 韩国车外观拉风 日间行车灯像两个大眉毛酷酷的！很适合做年轻夫妻的家庭代步车！【内饰】内饰一看就有一种不上档次的感觉 到还算大气！只是没换大屏之前控制面板全是红红的 看着不舒服！【性价比】性价比非常高！保养便宜 该有的基本功能都有 天窗 多功能方向盘 无钥匙进入 无钥匙启动！已经很满意了！但是后排没有空调口 不是真皮座椅 没有中控大屏还是让我有点小失望！【为什么最终选择这款车？】买车之前看了轩逸 宝来 卡罗拉…但是看到k3之后外观好看 动感 主要的是价格便宜 便宜 便宜！看到k3到把它买下来一共花了3个小时！【其他描述】不知道什么时候车门上已经有了一个小坑！是不是车漆软啊 门把手上的按键在洗完车后会失灵一会不知道是不是只有我的车这样！异响什么的问题还没遇到！|http://k.autohome.com.cn/spec/19724/view_1108077_1.html?st=95&piap=0 2886 0 0 2 0 0 0 0 0 1#20160510|2016-05-27
기타|2466656783|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 21:07:26|2016年05月15日 发表了口碑|来自：汽车之家Android版  2016年05月15日 发表了口碑  口碑    《十万左右性价比比较高的一款车了吧》             【最满意的一点】最满意的是后排的空间 后备箱的空间 还有我喜欢的黑色内饰。【最不满意的一点】买的自动挡的 动力比较弱 超车真的很费劲 还有k3的车漆 真的不敢恭维 小石子蹦都能蹦掉一大块漆 还有它的胎噪 不是一般的大 隔音也不咋地 还有就是后排座椅不能放倒 如果需要载比较多的东西的话会比较麻烦 不怎么实用 希望以后可以改改 比较是家庭用车 空间还是很重要的【空间】前排的空间还行吧 挺大的 但是后边中间有凸起的地方 做三个人中间那个肯定不舒服 【动力】自动挡的 动力比较弱 超车什么的一般般吧【操控】减震特别硬 起步的时候车头有异响 不知道怎么回事。十万元左右的没什么操控可言 都差不多吧【油耗】油耗还行吧 城乡结合部 7个油左右 在高速上5.1 也不知道油耗准不准 下次加油我清一下试试【舒适性】座椅怎么调都不舒服 一般吧 皮座椅是后加的 比较吻合 还打了气孔 【外观】韩国车卖的就是外观 k3k4k5都很好看啊【内饰】一般般吧 硬塑料的地方比较多 看起来很廉价 摸起来很硬 但是有我喜欢的黑内饰 这是我选择k3的主要原因之一【性价比】十万左右的一共就那几款 英朗 福睿斯 朗动 朗逸 起亚等等 k3的性价比偏高吧 适合上下班代步【为什么最终选择这款车？】看过英朗.福睿斯 卡罗拉 宝骏560 哈佛h6 本来就打算定福睿斯了 51和姐夫一起去车展看福睿斯的 姐夫说福睿斯不咋地 屁股太丑 16款的k3还不错 然后我就考虑了一下 就定了k3 因为价格都差不多 都是代步用的 所以就定了【其他描述】到现在跑了1300公里了 各方面都还可以 油耗也没有认真的算过 没了就加 缺点就是车漆真的很薄 伤不起啊 害得我只能去补补 但作为一款10万元左右的车型 k3还是比较满意的。|http://k.autohome.com.cn/spec/25737/view_1114009_1.html?st=77&piap=0 2886 0 0 2 0 0 0 0 0 1#20160515|2016-05-27
기타|2466656786|Autohome_review|K3(起亚K3)|ZHO|2016-05-27 21:07:26|2016年05月16日 发表了口碑|来自：汽车之家Android版  2016年05月16日 发表了口碑  口碑   《总体家用还可以 动力输出较为平顺 》   【最满意的一点】空间在同级车还算可以 主要外观好看【最不满意的一点】早晨异响严重【空间】空间较同级车我觉得还是可以的 唯独缺点就是后排不能放倒【动力】如果加速超车只要敢踩油门还是可以的 在市区加速较为平顺【操控】精准度还不错 就是方向盘握的地方比较低 有点够不到转向灯和雨刮器 过颠簸路段时基本还可以接受 后排过滤也还能说的过去【油耗】预期油耗在7个左右 不过一直在市区跑8个也还能接受【舒适性】座椅的舒适性还是满意的 后排还有杯架 【外观】外观是最满意的地方 因为够年轻 够时尚 符合年轻人【内饰】用料有点吝啬 基本都是硬塑料 只有门扶手是皮的 个人感觉在10万左右的合资车也还能接受 【性价比】基本还可以 在合资车算中上等了 家用肯定够了 性价比在同价位的合资车里个人觉得还不错 适合年轻人【为什么最终选择这款车？】买车的时候还看的丰田卡罗拉还有大众的浩纳最终选择k3 就是价位空间还有较为帅气的外形【其他描述】|http://k.autohome.com.cn/spec/19724/view_1114776_1.html?st=74&piap=0 2886 0 0 2 0 0 0 0 0 1#20160516|2016-05-27
기타|2466713280|Autohome_review|랑동(朗动)|ZHO|2016-05-27 21:41:02|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=180&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-27
기타|2466730834|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-27 21:52:01|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=218&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-27
기타|2466739629|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 21:58:02|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=122&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-27
기타|2466788773|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 22:29:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=185&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2466788952|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 22:29:02|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=116&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-27
기타|2466789283|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 22:29:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=167&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2466789396|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 22:29:02|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=123&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-27
기타|2466811444|Autohome_review|랑동(朗动)|ZHO|2016-05-27 22:43:03|2016年04月27日 发表了质量评价|"2016年04月27日 发表了质量评价  质量   该车主目前没有发现质量问题       2016年04月26日 发表了口碑  口碑    《朗于心 动于行》           【最满意的一点】当然是他的外观 流线型的身材 犀利大灯 日间行车灯 包括后视镜自动折叠 一键启动让人怎么看怎么喜欢 百看不厌 看了朋友的马三 b50|更加坚信还是咱滴小狼好看 油耗感觉特别省 非常满意 内饰比较符合咱小青年的眼光.（冲动是魔鬼！谁说的 朗动当前 把理智抛到脑后吧！）朗动广告宣传页上写的 我想说选择它不是冲动 而是深思熟虑过后做的选择【最不满意的一点】有点小异响 异响有时候有 有的时候又没有有点莫名其妙 胎噪 有点大 关上窗户 放点音乐还不错。悬挂我就不说了 广大车友都有体会 既然选择了它 就要接受它的缺点 哪有十全十美的 是吧！【空间】空间家庭用车应该够用 如果后排座椅能放到那就完美了 不过前排表现有点一般 反正我170的身高感觉挺好的0.0【动力】1.6自然吸气你还想和涡轮增压的或者排量高的比 不过1档有点肉 转速上去2档和其他档位提速挺好的 但是对于我来说够用了 咱开的是车 一个代步工具 不是灰机【操控】操控感觉不错 转向很明确 车速上来方向就会有点沉 为咱安全着想不是 喜欢他的油门踏板 踏上去很舒服 开朋友的英朗 感觉太抠了油门踏板做的一点点.还是小狼驾驶起来舒服【油耗】油耗特别省一直显示5.8|跑过一次长途来回900多里路 油才用了100多块钱 挺实惠的 天没亮出发 走到吃了一顿饭返回 头一次跑长途 还挺兴奋 小狼也给力安全返回 使我对他更有信心 更见让我相信选择了小狼我不后悔 油耗这方面非常满意【舒适性】舒适性方面挺满意的 腿部收放自如 感觉也不是很累挺放松 驾驶起来关上车窗声音挺小 开起音乐挺享受 真皮座椅舒适度正好 后排空间挺大 大家都说头等舱的感觉 【外观】外观这应该是大家都看好的一点吧!高大上的感觉 看大家改的前脸 后唇就是一部超跑在眼前啊 它腰身流线型的设计 耀眼的led日间行车灯 动感的轮毂不得不佩服现代的设计师【内饰】内饰.还是看中了小狼的炮筒仪表盘 以及做出了白外黑内的选择 特别突出的是它的剃须刀式的大中控台 布局合理 动感十足 包括整个中控台的用料以及设计非常喜欢|眼镜盒 遮阳板 正驾驶和副驾驶遮阳板都配备了一块小镜子 方便女性化妆 挺方便【性价比】相对而言朗动的性价比还是挺高的 可以和其他车比较一下 再者看它的销量就知道广大车友的选择是对的【其它描述】希望现代朗动配备全系ESP|紧急时刻保护安全的配置 相信以后现代朗动的销量会更好 对了最近现代推出了领动 做保养的时候刻意感受了下 配置 外观以及内饰的话我感觉还是自己的小狼更胜一筹 领动的内饰感觉太老套 都说车漆有点薄 这个没啥感觉 刚提车的时候碰过一只大羊 因为是新车不 后面还有跟着的车 不敢急刹 撞击力度感觉还挺大 除了前机盖有一点漆面脱 日间行车灯里面卡口松落没啥问题 去了4s店 维修人员给我免费维修了下如外检查了下外关 服务态度不要错 可见现代的车质量还是挺可靠的。【为什么最终选择这款车】当时比较的车还是不少 k3 朗逸 卡罗拉 英朗 科鲁兹 逸动 k3和朗动差不多 感觉还是喜欢朗动 朗动的外形 内饰 配置和性价比一直吸引着我 所以做出了正确的选择 选择了它【保养】前几天做了二保换了高端机油当时店里给我拿出几种机油我选择了一款中等价位的328元黑色的记不清是那个了没办法给大家分享 抱歉 还了油塞密封垫 空气滤芯 发动机机油滤清器总成 还有一个发动机润滑系统保护剂 正好有活动二维码抽到一个机油85折 以前活动领到的保养卷除去这些花了471元大洋 售后服务挺不错的 还给洗了车 不知道有没有被坑【缺点】A柱有点遮挡视线 车友们多多少少都有一点反应 转弯的时候大家尽量多注意下 毕竟为了大家的安全着想.还有一点 大灯晚上行车的时候感觉灯光不是太亮。"|http://k.autohome.com.cn/spec/20616/view_1089896_1.html?st=179&piap=0 2764 0 0 2 0 0 0 0 0 1#20160427|2016-05-27
其他媒体|2466812677|bitauto|易车 > 问答 > 问题分类|ZHO|2016-05-27 22:44:01|雷凌和k3哪个好|雷凌和k3哪个好     提问者：付建强  分类：  丰田  雷凌  买车  选车  浏览[5] 来自：易车手机客户端  2016-05-27 21:31  举报   雷凌和k3哪个好|http://ask.bitauto.com/detail/6599117/?leads_source=p029001|2016-05-27
기타|2466835339|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 22:58:01|2016年05月18日 发表了口碑|来自：手机汽车之家  2016年05月18日 发表了口碑  口碑   《热爱我的热爱 雪佛兰科鲁兹》   【最满意的一点】1。最满意的当然外观啦 当初买车就是看中这车外观成熟稳重。2。就是操控 对于我来说操控表现游刃有余。3。就是空间和舒适度 地盘偏硬 过弯悬架支撑到位 座椅软硬程度对我来说刚刚好。后排空间宽敞。【最不满意的一点】就是隔音效果不怎么好。至于油耗就是仁者见仁智者见智了。【空间】空间对我来说非常满意.【动力】我觉得还好、只有肉人没有肉车【操控】转向指哪打哪。我开着很有感觉【油耗】差不多【舒适性】就是高速噪音有点大【外观】相当满意【内饰】对于现在工艺水平就有点落后了【性价比】物美价廉【为什么最终选择这款车？】选车看过宝来 速腾。卡罗拉 k3 朗动。但是对比之后还是觉得小科适合我【其他描述】|http://k.autohome.com.cn/spec/14284/view_1122093_1.html?st=118&piap=0 657 0 0 2 0 0 0 0 0 1#20160518|2016-05-27
기타|2466835470|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 22:58:01|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=58&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-27
기타|2466881562|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 23:29:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=187&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2466881635|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-27 23:29:02|2016年05月24日 发表了口碑|来自：手机汽车之家  2016年05月24日 发表了口碑  口碑   《总体不错 一年跑这么多公里没被抛弃过！》   【最满意的一点】油耗 发动机 底盘！【最不满意的一点】变速箱挂档的时候有异响【空间】说大不大 说小不小 坐在后面一拳四指的空隙 本人身高1.78体重190.肚子像怀孕6个月的哈哈！【动力】一档有点跟喘不过气一样【操控】挂档顺畅 个在人开 没像论坛上说的有顿挫感 除非你换挡的时候离合没踩到位 不舍得给油门 毕竟是紧凑型车 不能跟大排量b级以上的车比 b级车以上的车能买紧凑型车一个半到很多！【油耗】高速夏天5.5百公里 市郊国道4.5不是吹的 市区7.5毕竟车轻了 但是多了esp 负车架用了全铝车架 发动机变成了全铝发动机 配件在升级 也算没简配！【舒适性】比老款舒适多了 最远18小时跑到贵州铜仁！【外观】苗条上的大气 大气上的苗条 尤其后屁股仔细去看性感中的闷骚嘿嘿！【内饰】就那几块破布 通用缺这点皮料啊 有点太抠了！【性价比】104000合资车的性价比不错了比大众厚道s【为什么最终选择这款车？】选这车之前看来过 大众思柯达 飞翔 日系车没考虑 现代k3 因为不喜欢大众的简配 飞翔的板车 现代的技术落后 最后去雪弗兰店想提创酷的 创酷的内饰叫我很失望 老爱唯欧的内饰！最后旁边停着一辆车 销售人员介绍过之后才知道克鲁兹新款的改进变化 直接订车 之前来过6年的的摩托 以前是摩托迷 后来换成车 微型车比亚迪f0 目前32900多公里除正常保养无问题 空调有时失灵希望以后能改掉 估计是通病！【其他描述】|http://k.autohome.com.cn/spec/19917/view_1129740_1.html?st=59&piap=0 657 0 0 2 0 0 0 0 0 1#20160524|2016-05-27
기타|2466884625|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 23:31:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=168&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-27
기타|2466884763|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-27 23:31:03|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=124&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-27
其他媒体|1602465885|zhidao_baidu|生活|ZHO|2015-01-09 04:16:01|东风悦达起亚k3是一链起动机的吗|我要回答分享到：|http://zhidao.baidu.com/question/1639094791051315180.html?entry=qb_browse_default|2015-01-09
其他媒体|1602807685|163|网易文化论坛-彩票大赢家|ZHO|2015-01-09 10:58:01|[好用]win7 64位 穿越火线[新版|"玩武魂延迟高用什么加速器  完美上线：穿越火线最新透视GG 2009年10月30日更新 每日更新 穿越火线最新透视GG 大飞 蜗牛 全部采用新算法 全部免费破解使用中。 下载地址： http://www.pk38.com/ color=#ff0000 size=4>本站的免费破解的穿越火线 好请帮忙宣传一下 不好请告诉全世界  【[好用]win7 64位 穿越火线[新版]win7 64位 穿越火线详细介绍】 版本号:v0.4.5|更新:修复SX错误|植入新的自动反TP功能.为了满足一些网友强烈要求所更新的最终版本!1.辅助功能键  F5地图透视|F6人物透视|F7准心|F8显鬼|F9人物上色|F10颜色透明.2.常见问题  游戏中按键无效的话|请退出游戏后重新尝试启动|或把  360保险箱和瑞星卡卡助手关闭掉.3.缺少文件 　　开启辅助程序后直接进入游戏即可! 　　游戏中按键: 　　F5地图透视|F6人物透视|F7准心|F8人物上色|F9颜色透明. 　　游戏中按键没反应的话|请把360保险箱和瑞星卡卡助手关闭掉. 　　缺少文件: ---- (有提示再操作) 　　如果出现缺少d3dx9_37.dll的话| 请运行大飞透视补丁 　　自动开枪（说明） 　　准心对准敌人自动开枪 暴头率增加75% 　　启动成功后 f7开启 暗黑3加速器f8关闭 进游戏之前需开启 否则进入游戏后快捷键无用。 　　如使用窗口化 请将桌面属性分辨率调整为1024*768 再配置自动开枪参数为1024*768  　　游戏里面无需设置 保持默认800*600。如不使用窗口化无需设置！ =============================================================================      【最好的[好用]win7 64位 穿越火线[新版]win7 64位 穿越火线】是由奇虎公司推出的完全免费的安全类上网辅助工具软件 它拥有查杀流行木马、清理恶评及系统插件 管理应用软件 卡巴斯基杀毒 系统实时保护 修复系统漏洞等数个强劲功能 同时还提供系统全面诊断 弹出插件免疫 清理使用痕迹以及系统还原等特定辅助功能 并且提供对系统的全面诊断报告 方便用户及时定位问题所在 真正为每一位用户提供全方位系统安全保护。点击下载穿越火线杀毒 　　穿越火线版 更新日志 　　新一代木马云查杀 　　-搭载新版穿越火线云查杀引擎 通杀活马； 　　-使用新的木马评估技术 更精确的识别和打击木马、病毒； 　　-安全专家潜心研制的木马特征识别技术 大幅提升侦测未知木马的能力； 　　-特有的威胁感知技术 能有效解决木马绕多传统扫描引擎侵害系统的问题； 　　软件管家 　　-优化开机加速：增加优化过的延迟启动与一键优化 　　驱动防火墙 　　-结合云查杀引擎 智能拦截恶意驱动加载 保证系统内核安全 　　漏洞补丁 　　-优化vista、win7补丁检测速度 　　-提升补丁升级成功率 　　本站提供穿越火线最新版下载。 　　蜀门onlie的问题 　　诊断平台: microsoft windows xp  service pack 2 　　ie版本: internet explorer v7.0.5730.13 build:75730 　　计算机物理内存:503.48mb - 当前可用内存:241.28mb 　　100 - 未知 - process: stormliv.exe [暴风影音媒体控制中心] - c:\program files\stormii\stormliv.exe 　　100 - 未知 - process: zssnp211.exe [zsmcsnap] - c:\windows\zssnp211.exe 　　100 - 未知 - process: domino.exe [] - c:\windows\domino.exe 　　100 - 未知 - process: ppsap.exe [ppstream 网络加速器] - c:\program files\ppstream\ppsap.exe 　　100 - 未知 - process: qq.exe [qq] - d:\qq2007\qq.exe 　　100 - 未知 - process: txplatform.exe [tm20052[好用]win7 64位 穿越火线[新版]win7 64位 穿越火线] - d:\qq2007\txplatform.exe 　　100 - 未知 - process: tipsextend.exe [tipsextend module] - c:\program files\thunder network\thunder\components\tips\tipsextend.exe 　　100 - 未知 - process: 穿越火线诊断工具.exe [] - c:\docume~1\admini~1\locals~1\temp\rar$ex00.203\穿越火线诊断工具.exe 　　r0 - 未知 - hklm\software\microsoft\internet explorer\main|start page=http://www.pk38.com/ 　　r0 - 未知 - hkcu\software\microsoft\internet explorer\main|start page=http://www.pk38.com/ 　　r0 - 未知 - hklm\software\microsoft\internet explorer\main|search page=http://www.pk38.com/ 　　路面水涟漪。安静烘托着细雨的瘦削 低头已是鞋湿衣冷。残风闻寒 周身的冰冷将血液里的悲伤唤醒 突然很讨厌盛夏的赤裸 暴露了太多裸露的肌肤。我紧裹着衣服 畏惧那天空飘过的白眼。我将手机耳机塞在耳朵里 也许是因为自卑着 我忽然很小气自己的。 　　眼泪不听话的分开过去 颤抖的双脚每走出一步 都会踩成结局。我回头看那些没雨水淹没的足迹 老天背叛着我的走开 一如既往的汇给我难过。过去的那些背影缩小在瞳孔里 远远的温度依旧是遗憾 我像躺在一样 在每个夜晚。都会蹲在一个从前没有风的角落。 西安高新区加速器催生科技小巨人"|http://bbs.sports.163.com/bbs/lottery/492382441.html|2015-01-09
其他媒体|1603831991|zhidao_baidu|生活|ZHO|2015-01-09 22:30:01|东风悦达起亚k3有带eps功能吗||http://zhidao.baidu.com/question/919721137236407859.html?entry=qb_browse_default|2015-01-09
其他媒体|1615231913|zhidao_baidu|生活|ZHO|2015-01-17 07:42:01|东风悦达起亚k33458型号多少钱||http://zhidao.baidu.com/question/1797376892724809467.html?entry=qb_browse_default|2015-01-17
其他社区|1636190570|360wenda|已解决|ZHO|2015-01-30 15:41:02|东风悦达起亚4s店可以自带机油吗|东风悦达起亚4s店应该是可以自带机油的 不过最好还是用4S店的专用机油比较好的。此回答由  官方管理员   推荐为最佳回答。 推广链接00x用微信扫描二维码分享至好友和朋友圈分享到：检举 -->答答好搜问答团队最勤劳最可爱的答答28分钟前下面是答答童鞋给您的小建议 您看靠谱吗？初来乍到 弄错了您不要生气哦(*^__^*)答答小贴士相关问题南京4s店东风悦达起亚k3要首付多少可以上路2014.06.01查看更多关于的问题 >>|http://wenda.so.com/q/1422598134701960|2015-01-30
其他媒体|1658546144|zhidao_baidu|电脑/网络 > 硬件 > 显示器|ZHO|2015-02-13 10:51:02|东风悦达起亚*k3显示屏无线连接怎么用|东风悦达起亚*k3显示屏无线连接怎么用7 分钟前登哥3336 分类：电脑外接设备|http://zhidao.baidu.com/question/2117007144381267747.html?entry=qb_browse_default|2015-02-13
其他社区|1662905618|360doc|最新文章|ZHO|2015-02-16 12:37:02|玄空相逢系列 玄空子老师资料汇编|"作者相关# X1 h2 ^' v' Z: d8 W·二气取象法9 h4 k"" w! d- k' m8 W| r·刘文德卦技二十法相逢是缘解析版- G0 x- D( Z$ K' u5 d  @' c·卦身# X  I: S9  9 o) K- w* \7 ?·卦序的应用# {9 m. q% R+ H: j"" D1 u·六爻理论集9 I' M- u  J2 {* B·浅谈“梅花易数”在股市中的运用; t4 F( u- E( @5 I·随口断9 D/ Q3 D3 ^- H·相逢是缘讲八卦3 R# [1 ~& D5 h| T/ I·六爻预测的多重思维- L' ?6 N5 w% c! o7 P"" J6 M"" V·玄空子《仙易俏梅花》之事态卦变法/ @7 B#  4 w! j. w# y) I( s: }·玄空子股市大盘预测研讨; b7 H. a- W! z- S! o·玄空子卦气流转法+ r6 @# J: c6 u) y·玄空子老师简论鬼爻持世. C- j"" N4 T1 F| M7 P4 G; k7 ~/ `. R·玄空子老师五行看性格  @$ d. n3 w% ?·玄空子爻位说象占例解5 P( b# @6 @| r6 B- F·增删与梅花断终生作者相关: h7 o& v4 F  w4 v8 u 3 {- y; @7 m+ ~4 y 本文由天机阁 www.tianjige .net 整理  更多内容尽在www.tianjige.net( R8 U. _: n! s | F5 a1 o6 w* V6 I) Z) r 　　相逢是缘 又名神仙姐姐。1988年生人 玄空子老师门下弟子之一 曾得老师的真传秘技《仙易随口断》、《二气俏梅花》等。8 ?6 z: \4 B) }# @- @) ^! Y& t6 n# r$ v% e0 E/ o- \9 u! D: D  O2 z  D- m; D$ e% J9 u1 C9 P& @  d( l0 K- G二气取象法9 f1 C- ?3 H6 Y) o   N. U# X6 U4 i$ O' j6 A( j4 \! U5 Q8 O& g) k| [| n5 i1 \  X"" _  `7 R相逢是缘) K' D6 J( J4 b. j) @) L3 l) S7 K8 N) D$ m: @1 N* Q' G| K* e　　二气俏梅花是一种只取阴阳二种卦变 按1、3、5、7、9、11为阳 2、4、6、8、10、12为阴 通过笔划、数字、事物之阴阳 直接分辩出要测事物的阴阳属性 以简单至易的断卦方法 直断判断吉凶的方法。2 [3 a! ^8 q- {2 @$ Y5 w1 v| D+ F$ `| n  [( f　　传统梅花取体用。二气梅花可取可不取。但其易理至易至简。一般地 一般即出 以八宫卦分出其阴阳大气 然后再根据具体卦象进行分析。在实战中 实现化象具形 化形具义 直简断占。$ e6 y"" l1 w"" u0 W9 W+ d; `( a; T8 M9 c4 \- `; y/ U  e& V+ _- u. _6 z& _　　在五行取法上 有别于传统梅易 有以下数字。; [- `8 N4 ]# U- B5 ~  O"" e6 Y7 X# t"" s- q+ H3 v　　1、2为水。1是静水 地下水 2是动水 江湖河流。遇火成天上水 雪、雨、霜、雾。| j0 x2 t8 S! b- s( Q% v8 @/ E$ M- q! h/ G. b6 R' }　　3、6、9、12为土。3是大地土 6是墙上土 9是丘陵土、12是坟地坑地土。' i& z5 [3 _0 m2 a| N2 _: j4 H| D# x1 t)  4 c) @　　4、5是木 4是阳林木、木制家具、大树 5是阴木、花草、小树。! L0 C. }0 @+ K6 t$ `$ s1 v9 C6 U+ a( a/ @: f　　7、8为火 7是外火、太阳火 8是内火、7克力大 8克力小 如7克11力大 很危险。/ E1 W6 d. y6 {5 `$ F7 S. G1 `3 d; F# H: g5 P% c1 V$ _9 d3 c　　10、11为金 10为阳金 11为阴金。. N! `6 l2 Y- [$ Q/ J* l- O9 I"" ?& z* N+ @　　因此法我师还在研究阶段 还没有成熟 因此 不便全盘公开。而且 说句心里话 除个别基础好的 别人看了也暂时学不会 至少会学不到其精妙处。但有一点 梅易的取象法 在各派梅花技法中 是可以通用的。传统的 包括黄见的梅花 因其取象法的单一 不能详以至用 所以 一般的学者 若非有高深的功底 在占断时 有时并不能直接断准其事。; {3 r7 L3 `) z|  7 B2 J( h"" }5 t8 ^% O8 `4 {* s　　二气梅花将气象数进行了细化 细到了生活中 所以 在取象占断上 是有别于其它的。并且 这一取象法 完全可以为它法所用。# ^"" r( ~% [| Z  t3 J"" }.  * K4 Z7 e3 \- P1 u　　我今天主讲的取象法 是空象的取法。关于空 大家在六十甲子中 在六爻中 都有过应用 旬空 月破 非常至简。实际上 梅易也有空破。如果象一些人哪样哗众取宠 也来个《梅花新大陆》 那么 我觉得 我老师的这一取象法 也称得上是新大陆了。; q0 f( y8 ~) }4 ?"" b/ p2 z3 h0 n| S& z' e3 k　　关于空破 在梅花中怎么取？非常简单。以今天为例（癸丑日） 今天是寅卯空 那么 卦中出现震、巽卦 就是空。破我不用讲了吧。本月中卯木破 对应就是 巽为破。知道了空 有什么用呢？大家知道 金空则鸣。木空则朽。土空则陷。火空则升。水空则流。在一个卦中 体卦出现了空。结合实际情况 可理解为 他心里发空 不在本地。测工作临空 是失了工作。测官运 官让人家得去了。然后结合我前边提的五行空法之用。金空大发雷庭。土空痛痛苦不堪 无力自拨。由空象 可看出许多故事。如果你看到木空 在给一个人看卦时 可断为 坏了心肠。腹中无物却目中无人。因木是离火目之原神。水空则是他要走 工作的变动 逼走了他。这里 我们在断卦时 就有了更多的象 在占断时 就会更生动。& V6 p| f0 G7  . z$ U| b7 n2 P; ?- x"" s* Y4 d　　一占例讲解。 乙酉月　乙酉日 （午未空） 地风升　　　　 雷泽归妹 　　　地天泰　　　　 　▅▅　▅▅　　▅▅　▅▅　▅▅　▅▅　 ▅▅　▅▅　　▅▅　▅▅　▅▅　▅▅　 　▅▅　▅▅　　▅▅▅▅▅　▅▅　▅▅　 　▅▅▅▅▅　　▅▅　▅▅　▅▅▅▅▅　 　▅▅▅▅▅　　▅▅▅▅▅　▅▅▅▅▅　 　▅▅　▅▅　×▅▅▅▅▅　▅▅▅▅▅: K  x1 ~' x% i3 _5 A  \! x| Z/ X　　这个卦 是我老师给我讲解时 举的他的一个占例。这是占婚姻的卦 是他所在地方 电视台的一个记者 通过他的妻子找到玄师 在电话里 我老师按当时的时间：4.05随机取出此卦。老师的妻子 也是一个记者。; E! p& Q2 a| Q. B| l$ Y) H! L  ~3 {7 L1 D1 w% R8 ?　　断：现在你的女友不在家 不跟你了。; a2 Z; e) r| P5 Y; g: V% X. _9 b) R"" M) N- h! v　　乙酉日 寅卯空 本卦中 坤土为体 巽木为用 为他的女友 临空。# A( h3 z  L) X+ q! R3 A"" N0 S| Q& }3 x  V( q& H　　为什么不跟了？而不是暂时出差或回了娘家？日月双克巽木 动又化回头克 这是有去无回。$ O( [9 N| c8 A"" a* `"" ?8 e/ E* u"" f　　那为啥不是死 而是跟了别人？巽木临空 不受其克 只是不在跟前 空者 她在这儿是受克 她跑一边去了 不受克 所以 没死。8 z$ o| L9 o+ ^& d# g$ m/ L) ]8 k8 _& a7 y; L/ i| j　　这一点 大家理解了么？打个简单的比方：  _) p; E& q5 M: c' f| s8 m; S"" O4 n"" j* S5 p　　插：就像六爻的旬空避克。4 p8 [) [6 e& E; O: \$ z6 c: }# t3 W　　对！伊拉克战火纷纷 人在那儿 说不定就死了 可这个人跑中国来了 到这里听来了 所以 没事 但在伊地 还是克重。换言之 如果他不空 就完了 必会克死他 而且 这里还有一个大家要知道的 互卦有震木相助 用卦又动。动后怎么样了？地天泰 她跟别人泰去了。( `| _: a( D% i1 x4 A$ W5 B1  / f7 o　　当时 卦主问我老师 你说：我与她成过几次 分过几次？这个几次 怎么断呢？巽木克坤 坤是卦主 为负三数 断 三次了。+ w' X/ q6 O| G; u) f. b; m4 C- v$ _% J) ^| i( b　　巽木之互为兑 克巽为其官 兑为小 第一次 因为钱 巽木克土 土为巽之财。体互为震 为夺财 震为长男 你哥哥跟你借钱 你女友不高兴了 离开了你。大家可能问 为什么这是第一次？ 因坤为母 代表万物之始 所以是第一次。. W7 k' `  a9 y% C/ u6 ^* B# W& v2 k( P; [: ?　　第二次 下互兑为二 下互 也是接近之意 所以 取为第二次 兑金为克巽木者 为其夫 所以 第二次是跟一个小她的男友走了。卦主答：是的 他们在一起后 经常加架 我劝她 她又回来了。. U( ?2 d| U  ]3 d2 V9 @9 n. i9 X　　问：第三次呢？跟一个有钱人走掉了吗？呵呵！* \' [. g| ^2 ~$ ?. P! o2 P3 P( h. m7 f　　答：对。第三次 不用我说 大家已经看出来了 就是变卦之乾 这是个官 但他在坤下 我说了 坤是用卦之财 他生乾 所以 此人是生意中有钱 是企业老板。) f3 E) T"" f- s| `# q% _1 o5 n$ Z4 m　　虽然大家都知空破 但是 不点破窗户纸 可能许多梅花易友并不知道空可以这么用。4 S0 M$ n& V4 i*  ! Z"" s2 I$ r$ U8 ]6 q8 r# l( c$ \. K) J5 F　　问：有一个人 此时是得肝病 现在正在病危 在手术台上 那可不可以救的回来呢？（若是以今天讲的课为基础的话 以这个理论来推。）5 M2 {# z8 B5 o7 n1 ~% C6 t7 P  p' H　　时间：乙酉月　乙酉日 起挂得火雷噬啃 变山雷颐  火雷噬嗑　　水山蹇　　　山雷颐 　 ---离火　-　-坎水　---艮土 [用]-　-　　　---　　　-　-　　 　 ---　　　-　-　　　-　-　　 　 -　-震木　---艮土　-　-震木 [体]-　-　　　-　-　　　-　-　　 　 ---　　　-　-　　　---& C- T2 O( Q| B- j"" U"" K. L4 j4 c% [* _; X8 }1 s　　这要结合具体情况占断 如果看此 我看此人 没救也。震木被日月所克 病很重了 互中有坎水 是靠点滴维持（是 在手术台上 大量输液）。上离火 现在神智不是很清（嗯 重度昏迷） 上互坎水 下互艮为山 变卦山下埋震木  不用我解释了吧。/ m2 ^: i9 E# a  o/ m$ ?$ P4 R2 Q( P| k5 K8 P! C9 M! \| C　　插：山雷颐------好像一口棺材。& M+ l$ l6 {$ d1 t1 K4 u9 z# n"" u. v& m  M0 h　　答：对的。/ F"" R| M( R+ n7 v5 ?: D7 I| Y! s"" c| b7 w# q% k3 H　　问：若是变为震为雷 是不是还有一线生机？但此时是空亡 那是不是也是没救呢？$ i! R3 O9 M7 F8 S9 e5 _- I- a7 E  n8 b8 K/ v/ o6 w　　答：变震就会没事了。2 P1 a1 ~| a& a9 j4 F( D2 m4 i| z. e* u- b+ s8 u& k2 L: R2 q% Y　　问：大病为空 为退去 加上变卦比合 所以为吉吗？9 {6 }; J* b) o4 w) L% Q4 t2 `6 ?: i0  8 K3 a. _( ]- y8 }0 G　　答：可以这样理解 但很久起不了床 只是 没有这个假设 你给我的卦 变是这个。刘文德卦技二十法相逢是缘解析版' H8  8 M* o/ Y1 f$ F$ [7 P: l' j) ^   m. l1 b2 H( N7 ^"" @0 _/ f % q& J9 }7 V8 ^& A8 c 原著　刘文德 ! _! F2 [5 O6 D! A( C! a% ?/ Z4 n) \& n4 u| m/ L解析　相逢是缘 整理　小飞熊( E! \  C  K$ m8 I6 `"" a' G7 g  L' _( l8 x二00七年三月八日;  / K: F# ]8 x1 q8 j: b6 Q8 K9 ]"" h4 D! Z8 T9 p' H　　刘文德的卦技二十法对于六爻学者来说 具有较高的学习价值 是提高六爻预测技艺必不可少的技法之一 但因原文中诸多地方不易理解 相逢在自己的群中 进行了讲课试的解析 将陆续传给易友把玩 转贴请注明出处。0 }( o0 j/ N| E! W; M- t$ ]$ w) [& ?5 u' Q　　一、场态观卦4 `: @) O$ D! k8 Q7 b) v6 A: ?5 k7 X　　什么是场？场就是环境。人有生活的环境 卦有生存的环境。一个卦所在的宫为大环境 大环境是一个虚指的概念 如经济环境 生活环境等 但它又是无所不在的 引领卦的气运。上下卦为小环境 小环境是一个家 一个具体的场所。你做生意 整个大的经济环境不好 你所在的市场 也会受到影响。影响力的大小 卦中看 就是日月四时的力量。小场制约三个爻。三个爻 因为我们常看的是用神 同宫中的其它爻 它与用神的关系是 他们是用神的邻居。而另一个卦中的其它爻 如 用神在四爻位 三爻位的也是邻居 但这个邻居同一个楼 另一个单元的它与用神所在的小卦的另外两个爻不同。9 N% A/ F9 [; f. a| G6 C| @! \* c　　尤其我们测比赛类 对这一理论能更好地理解。世应是双方。他们不可能在同一个经卦中 那么 他们所得到的力量就会有所不同。我们习惯的看法 是先咬用神。有了场态的观念 就不同了。因为“场”对爻具有一种作用力 所以观察“场”的时候 把时(年月)、空(卦的环境)联系起来看 各种作用力的表达就会更清楚了。一个人在国务院工作 又逢盛世 那么 他就算是一个普通的职工 他说句话 也非常好使。把不逢时的皇帝放在监狱中 他就是平民一个。由此 我们知道了 一个卦爻 不只是日月对它有益他才具有较强的作用。如果环境不是很好。也会使他的能力难以正常发挥。一个人 上级任命他为本县的县长 他在这个县里 非常管用。他到海上的轮船上去指挥船员 可是他的话只能是屁话 没人听他的 而他身份没有变 他还是县长。- T8 m5 ~| h! m6 j; U6 L. O) l) X' g+ w- {* m| a& d9 s6 M# ?| t| X　　例：八月问官职及调动情况得“地雷复”之“地泽临”；酉月 8 Y6 I( b% O  Y3 e& o$ {6 j# G; ?- M  @| ?7 j. f; t　　　　　　　 地雷复　　　　　地泽临 　　　9 W: t1 V4 B+ v3 n7 Z! x3  8 @- q! d. }　　　　　　　青龙 子孙酉金 ∥ 　　子孙酉金 ∥ 　 　　　) i! m- w. q* ~; I) X( S0 Z% g5 }0 L. O6 t| F' \% c; W% A　　　　　　　玄武 妻财癸亥 ∥ 　　妻财癸亥 ∥ 应 　　　# w2 _1 @4 G9 g# w& {2 V5 x2 r7 N"" `- j4 D7 D　　　　　　　白虎 兄弟丑土 ∥ 应　兄弟丑土 ∥ 　 　　　: ~3 f' ^( D8 f( x9 O9 f4 J8 R8 P9 G"" w: \　　　　　　　腾蛇 兄弟辰土 ∥ 　　兄弟丑土 ∥3 P: ?"" _7 Q1 Z+ ~+ f- ^& \8 _& f! J& C"" z　　父母乙巳：勾陈 官鬼寅木 × ! ]( R8 H7 A6 r& l: v* N0 C0 v4 J"" K' h"" r# B& C- }* X$ A( t2 E　　　　　　　官鬼 卯木 ／ 世 　　　& y: a"" H: H5 T# q5 n0 y+ R# z) w* c) v( O/ y　　　　　　　朱雀 妻财子水 ／ 世　父母巳火 ／0 S5 r"" G$ b& T/ q# n"" }$ B0 @+ u"" l' W3 T- }+ @6 e) N　　刘文德原断：用神官寅在震宫 这位先生在本单位 职务还是颇相称的。但“震”卦这个“小场”被月令所克 目下单位不景气 连向职工发工资都常从外单位告借而维持（外卦亥水的财来生合内卦的寅木）且常有口舌是非（震为吵 兑为口舌） 震变为兑 调离本单位后 虽然能在职务上升一级（寅变进神卯 卯又是正神） 但变卦后 兑金克卯木 故必将在新单位中受挫。兑为女人 为口舌 比皆为受挫之由；加之变卦兑金的场克卯木的作用 故入新单位后好景不长 很快处于无实权之状态。5 d! E9 A: `  B"" e% U: R6 m' c. L5 }) T2 ]# b( p　　原断中 我们思考以下几个问题。# \& k. e/ A; U2 V; N7 h"" k8 y. E"" X3 @1 T&  　　1、 变卦的卦宫 能够对原卦产生影响。9 A  ~9 T) T1 V$ o# i# J. `/ c7 _6 c! b. X3 K* p1 P　　2、爻的变爻 是事主现在时的延续。而且 动必有因 它也是事情将要发生情况的指引。 由此我们知道了 动爻 往往是破解卦的不吉 解灾的重要地方。就是说 他要工作动 才会有没实权的待遇。如果他不动了 就不会有了。非常简单直观的解灾。 　　3、变爻是末来时 它在一定意义上讲 它所指引的方向 是对末来的一种指引。 4、工作场所 我们常用的方法是 以应爻为场所 以父爻为单位或所在的场所 在实际运用中 所在的卦宫 就是场所。第一例讲完。 　　　　　　　　　　　: k5 ]+ R! Q* A/ r0 _9 O% q3 s' i6 s7 W( u$ R| ^% r　　二、卦象拓扑/ P; U5 O1 y0 c* Y' M' j7 x+ Q; W% d9 v7 Z  u2 K　　拓扑 就是把卦改变形状 再看它象什么。一根水管 你把它从中间割开 它的构成的本质并没有改变 但是 形状变了 这就是拓扑。| e5 J4 g0 Q8 n1 k3 Q- r+ W0 l4 O1 V　　比如震卦 震为车 是因为 你把底下的一阳当成了地平线。上边的两个阴爻 象四个轮子。所以 成车形。在断卦时 特定的情况下 我把震看到水池 也是此理。下边的一阳为池底 上边的阴爻就是水。同样的卦 只要我们善于联想 结合时空一个卦可以拓象成许多东西 震为气体 气一般由水而来。一阳初升方为震 是阴气至极后阳气的开始 所以 把震看成水 有它特定的卦象意义。4 E2 X  x5 h% C# v: E9 H. g' ]6 @! R8 }' ^! H; r! ?　　当然 卦的说变化要合乎法度 方为卦理: z  Z! ^6 W8 i% n)  : A8 K7 \7 N5 q　　例：壬申年巳月癸卯日申时 一妇问遗失100元之事。起“蹇”之“谦”$ f5 \"" K( h' g  {% b* C; `$ g& G# W! y% W! y1 @"" J5 T$ a　　　　　　　水山蹇　　　　　地山谦# A& z7 n2 T- K2 f; T"" P$ C"" n% @; ?% i# c4  7 J　　　　　　　白虎 子孙子水 ∥ 　　兄弟酉金 ∥) s) Z' a9 t6 K: h$ d# @"" X* g8 U"" O9 g7 n　　　　　　　腾蛇 父母戌土 ○ 　　子孙癸亥 ∥ 世0 ~% i( G5 d$ k4 k/ N% X. I  @| P"" r　　　　　　　勾陈 兄弟戊申 ∥ 世　父母丑土 ∥7 Z  ?: d5 D5 a: i( d$ m| m. H. u( Y% V% @+ w3 C　　　　　　　朱雀 兄弟申金 ／ 　　兄弟申金 ／2 }+ W5 W. e2 P5 x. w8 m| V"" V- d2 ^6 {0 s  _　　妻财卯木：青龙 官鬼午火 ∥ 　　官鬼午火 ∥ 应6 D9 N' A* P- e* r0 U3 s9 m| N' t! a1 [  u# q; i　　　　　　　玄武 父母辰土 ∥ 应　父母辰土 ∥5 P0 b$ H1 I. H5 K*  5 Z3 x% _$ U"" h8 z　　1、财为用神 伏官下。; n  A) S! S% ~5 L. O5 h! q9 [: T| l/ t1 t2 B: `3 P* P　　2、官没动 而且此官临午 得日月双助 是光明正大的象 断不是贼人所为。) ~$ w| X( ~. C. q0 C5 r+ h| {4 p' f"" ?# p! G　　那么 此官就具备了另外的意义。财伏不动在内卦。二爻位为家宅 所以 此财没出屋。当天是卯日。引财而出 动爻来合。所以当天可见。) e"" H% @+ s+ y  r! J4 O) s8 V' @+ E% c$ i7 q2 e　　3、动变亥水。与财又是半合局 变卦所指引的 往往是时间的定量。所以 断为亥时会出来。8 H"" H. z"" _6 M5 \3 Z2 Y| i+ E+ {9 U6 \. _　　4、在什么地方呢。内卦为艮 是裤子的象。二爻是宅位 裤子的家是什么地方？裤子的口袋。这是把卦放大的看象法 由此 我们知道了 巽是裤头 兑是老头衫等等。象就出来了9 }. k| j+ o) i1 s- A9 k  c: t6 S3 g* U"" X/ Y  B5 B) }| p. V8 M2 X　　艮又为床象 为什么不断在床下呢？因为二爻不是床位。- D7 h6 ^1 M: O; ^1 Y2 `9 I4 U1 h& g% _　　一般地 在无其它爻配合的情况下 三爻为木才能定为床。其它的 都不能肯定3 w! j| V* r+ R( Y2 _9 C| S% e$ b* o8 l| q　　例：一个占得未济之损问职业$ u5 ?4 C: v% J"" @  C5 r0 P: t. `* G! c$ A' ]+ {　　　　　　　火水未济　　　　山泽损; T5 f: C/ L7 P; j/ p# X: ]! F2 n0 Y2 J; o! j7 A9 V　　　　　　　白虎 兄弟巳火 ／ 应　父母寅木 ／ 应' @1 T. F3 h1 c$ j. y; F5 L| ]2 l6 `1 a5 @: I& m$  ! J4 T2 A/ [( V0 J& `　　　　　　　腾蛇 子孙未土 ∥ 　　官鬼子水 ∥; G7 E+ q; H! Y: m4 d# N0 w( X& t6 ^- y% b' s( o& R' Z　　　　　　　勾陈 妻财己酉 ○ 　　子孙丙戌 ∥* Q) i+ W2 A' @"" Y$ `% v. v| R| z; M| m7 [# H8 r2 h: i　　官鬼亥水：朱雀 兄弟午火 ∥ 世　子孙丑土 ∥ 世/ a0 w1 k1 J: C; p"" v8 b"" C| M- m. h4 \1 \| A+ O+ ^6 A　　　　　　　青龙 子孙辰土 ／ 　　父母卯木 ／3 t# j3 m0  + L; o3 s$ Q5 Z8 b% j! X2 Q% s$ O1 e9 Z　　　　　　　玄武 父母寅木 × 　　兄弟巳火 ／- i  ]* [3 l# ]) B- p+ p5 z# U* J8 v9 o- G; I0 }9 \　　刘文德原解：此卦财临己酉大驿土发动 内卦坎为轮 父爻（车）动 说明在路上开车赚钱。开什么车？外卦（*图）形状象“拐的”（三轮摩托）的俯视图 所以此人是开“拐的”赚钱的司机( R' y# a| Q1 c! i5 b* r* a# Z0 o6 P# S0 n/ y　　相逢解析：3 h$ ?$ b  l4 t- s' X+ M* C2 Z7 F7 l& z/ v- r; S: u  `; a　　1、此卦原卦断得迁强。有后加工之嫌。"" Q& d"" _; Q) ?2 U) R| e| s8 K% s. G$ x5 @7 a　　2、父动化巳。动出之火与本卦没发生关系。那么 它有能力与主卦中的其它爻发生关系。查卦爻 正好与财酉有关系 此父即是财的长生地 又与之相刑。父代表车。说明什么呢。这个车 能给他带来财 也是个破车 老让他破费。9 e* q0 ]| ]) L3 }' J| f1 d2 u/ U& s7 j( p　　3、父在初爻临玄武。也主此车没牌子 是个偷着跑的车  B2 p( [$ g$ H) a! T' h% Z/ o% B$ o| p( k0 }/ i% B7 z　　4、五爻为正路 它动出之兄生五爻 而主象父克五爻 说明它不敢正经的上大路 而财与五爻这个路 贴身泄五爻之气 五爻被动地生财。说明是路上财。( W"" b% P2 y1 ]; f2 ^; g| q2 k/ Q| C$ i  {% _7 ^　　由此断定 此人的职业与交通有关系。( f4 R: u. Y% V4 @8 u) z5 s/ G8 O; T( m* P' T) _# _　　5、但车怎么看呢  a$ G) V' T1 l' x+ P: n6 K7 k""  ! J　　我在仙女群中讲过 一个卦是打开的太极图。它原本是园形的。那么 上爻就是初爻的邻爻。上爻 初爻 二爻 与代表车的父要构成离火卦。主卦加上变卦 两个卦其实也还是园形的。离为三。坎为轮。主卦的内卦就是轮。外互又是一个轮。初 上 五爻加在一起 还是一个轮 是三轮。- G"" U' {1 y+ U. V0 M: ]; q: B# {+ u. P$ w% I　　6、如果单按刘文德的那种化象法 说心里话 如果不是事先知道答案 我断不出来。) [! i  _4 T1 m) ^( @& r' ?2 ^1 Z+ f7 P% O- L; u3 o9 L$ ]! ^　　我不敢把财在离宫 就定为是开三轮车的 财动离变艮。也没看出车象来。6 j) U; X/ q% ?8 K| v. U| H- e& S2 o: o4 Z) e- B　　有了父爻是财的长生地这个前提 再结合其它象断 我才能初步看出一些门道来3 V! H% Z: T; n  f# u$ }2 x+ O' N"" M' R6 L; R4 }+ D| I　　例：癸酉年庚申月辛酉日 解先生求测家事 得鼎之小过。"" v0 J0 @: @( j1 C& w; A1 n/ y0 J8 E; s& d　　　　　　　火风鼎　　　　　雷山小过( ~& u  l  w1 e/ T3 h2 C# G-  / S"" N2 z(  2 T　　　　　　　腾蛇 兄弟巳火 ○ 　　子孙戌土 ∥9 f8 H; ]| L( m' H& e9 `! Z4 J# @9 z5 l9 w　　　　　　　勾陈 子孙未土 ∥ 应　妻财申金 ∥' l2 z* Z#  | }: E) ^$ p5 g4 a3 f5 c( S　　　　　　　朱雀 妻财己酉 ／ 　　兄弟庚午 ／ 世% j0 ^| {( w( ?/ R* H% k. J2 \$ O. Y( e　　　　　　　青龙 妻财酉金 ／ 　　妻财申金 ／. ]7 T$ i3 F' s% I| D1 r; a6 V& M$ d4 k: O9 a　　　　　　　玄武 官鬼亥水 ○ 世　兄弟午火 ∥. T# S* ]/ b; T8 {: {- [8 ]+ v% d# ]5 v7 L0 q　　父母卯木：白虎 子孙丑土 ∥ 　　子孙辰土 ∥ 应+ M2 S( B4 y! J| H8 B# o+ v3 B' O1 l; y  x) c! G! u　　1、断家事一般以世爻 财爻为用神。兼看宅爻。) X$ e' A& ]9 T9 t% q| }) ?- f$ k2 V/ J0 L2 }! v1 T+ O　　刘文德在断了此人家的一些事后。重点断了他家丢了一台洗衣机。: h1 U! d+ t% k| `& ?9 e9 D! o9 m. }; F: i: Z! Z% d| o　　首先 玄武临宅动化兄 二爻为家中的路。: A1 M) l+ L/ E' i"" l5 P$ S; x: f1 Z: ^6 j　　说明是在家中发生了与玄武和鬼相关的事。"" d; N' `' o. B. H& b- N0 _+ B/ W7  . b- i5 @3 Q　　此卦官爻持世临旺无伤。说明非伤灾类事。6 }"" B+ V# o5 }) L( h% b% l/ U  D  @| v6 k3 M　　那么 他求测的是家事 所以 也非工作类事。围绕家中的事展开。( K' n  P8 ]1 Z$ }| K  `6 D| N( l$ T  ]"" A2 q1 R( l7 E) u　　2、官代表死人或官司、盗窃。| q2 z"" b7 M( P% F( w! s$ r# Z# ^$ ]8 g"" d& ^% {- l- Z　　用排除法 我们知道了 官不受克 一个家中 也不会把死人放在屋里。所以 排除。而官司呢 是应该与应爻发生关系。应不动 不来克 世动化兄又与应合 也不应该是官司事。那么 兄鬼动 兄是劫财之神 他们合在一起 最大的象征就是盗窃。5 P6 H. @$ r  V+ p3 h"" V"" V"" ]* p* ]9 X6 ~+ D6 P　　3、丢了什么 在没确定是财或其它什么东西前 看鬼位不失为一个好的取象法。巽木的形状 打开来 象个小脚的橱柜。小脚办公桌 冰箱 都具此象。暂时还不能定为洗衣机。| T( g- ^/ `; R8 t"" b; G  j2 ~/ ?+ X6 Y5 y  t　　但鬼爻是亥水 水动了 水在柜中。亥字是个扭曲的象 如同衣服在里面搅。但这 我们还不敢肯定是洗衣机。结合梅花法。巽木为软 有衣物象。巽为风 变动后成艮 为止住了 止住后呢。亥水成了午火 干了。好比是洗衣机洗完衣服 甩干 停止以后 衣服就差不多干了; y& C+ x: ]: u3 J3 i4 V' U' G2 X9  % W　　这样一看 就把洗衣机的象 更清楚地看了出来。5  6 q) u0 W% p/ s8 y. O| ^: t( ]4 C   8 ]3 }% p0 y0  & S　　思考：- p| j(  "" U1 N# ]  A  \6 q& J5 F+ f2 S7 `( ?. _| r- d7 h2 X　　1、卦象的坤或乾 在高明的卦师眼里 是活的。它们在代表本身卦象的时候 还具有其它多种变象。6 ^. Q( M7 s- j/ ~$ E# B$ O' x3 k+ ~( D8 g""  4 H　　2、要学会从生活中现实象的角度去看放大 变形卦象。7 r& F  E0 m3 u/ n+ }"" n2 i! e% H9 l　　3、拓扑的放大与改变 不能仅就一个卦象去改变它 必须与其它的爻象、六亲、六神 甚至纳音等结合起来 否则就是乱变。' x8 X' F% H! T$ T6  : s3 m; ~3 O  b4 t  f0 ^7 D　　三、事态顺序. j9 Y0 Z8 t; b$ E7 X8 `6 H; g0 s3 K& {& G* g1 T! E7 }0 T% Q　　“大小运限 从初世起 阳顺阴逆 六位周流。9 U  B  Z6 [& P"" v# x% m% _7 q' S! J# Z; y) E5 H/ ?　　《易隐》-对于运限：“从正卦世爻 一年一位 在阴阳逆行之以定吉。阳世为顺 阴世为逆是指。一卦30年。一爻为五年。' O| Z3 @| L' `"" e3 X"" Q2 _) O6 Q8 x' a7 e| N& E7 e. e5 B! N　　阳顺则自世而上 阴逆则自世而下。 由此可知 事物发展过程可以把初爻作为事物之始 以六爻 为终。周流观看卦是一个园。上爻的上边 是初爻。; s& I2 k- m# M) O( Q# m/ V7 m6 z+ m; R  K! X　　1、假如一个卦 世爻在上 应爻在下 阳世 事物自下而上地进行 那么此卦反映的事端便是由应方先开始$ ~+ m( z5 k3 n% v9 u% Q% }; M; u( M　　2、阳爻表示过去 阴爻表示未来/ t1 t: J6 w7 m4 l/ _+ H4 N6 G/ a% j# A　　阴爻为阴性的 内在的 或暗昧的事 阳爻表示快速进行的事 以此为序展开。& `; p"" X9 Y3 n) ?0 R- A  q! k0 l1 h: Z　　3、事物从上往下进行时 有关卦象方面应当倒过来看' e; N' ^# Y$ ]) u8 }+ C$ u- i6 @% x: E6 A1 \) [　　4、在事物发展中 哪个爻发动 哪爻就有情况变化 % j4 Y' _+ A6 d3 z+ V2 _| O& {* i"" R2 l"" F　　例：癸酉年戊午月乙丑日 湖北某村一男人神秘失踪。3 N5 j* ]6 W' V6 m# \! y* v( h; i9 n4 _( ?2 r　　泽水困　　　　　雷地豫& V% U$ W8 Z* [7 R: a8 z7  4 U3 v' Q3 ^: E5 e1 L　　玄武 父母未土 ∥ 　　父母戌土 ∥2 P8 G# X% F3 n% J4 ^* V3 e% S2 _- o! c0 e4 U+ C- R　　白虎 兄弟酉金 ○ 　　兄弟申金 ∥% `4 A: s| t! p' {4 \7 d"" z9 K5 ?: Q6 _"" l3 @9 V8 z　　腾蛇 子孙丁亥 ／ 应　官鬼庚午 ／ 应| i( f! S# J5 L! K6 f# K- R% }3 _% q; N+ V$ Y& X# S/ {　　勾陈 官鬼午火 ∥ 　　妻财卯木 ∥/ Z& T* @. A0 B) u) B"" ^6    S  Y6 n  B; D/ z　　朱雀 父母辰土 ○ 　　官鬼乙巳 ∥* H0 C$ q( Z: a$ f2 K0 [$ ^  F; V7 X* T| K3 _& s. G　　青龙 妻财寅木 ∥ 世　父母未土 ∥ 世- Q5 @9 U+ W+ S$ m% T8 _( F% E| N. x: e3  4 d4 `　　刘文德原解：酉为门户 白虎临门户动 巳伏伤人之兆 此卦世爻为阴 故事态线自上而下。) b! p' q4 r3  $ n+ N4 m+ g3 P. G+ J　　兑为口舌 应爻空亡 玄武为始作俑者 故此人在家中与老婆呕气 老婆出走为事端为始无疑。3 x& C. N& K) O% K: a3 U4 ?* Z. X4 ~| B& o| b　　相逢解析：刘文德此卦解得不明白。9 t"" X8 J0 {6 `! Q) i4 a8 z9 c# W4 Y4 i& E/ G' M2 ]' c　　一是他怎么就看出是他妻子与他吵而不是别人？9 p% g) T| L. t8 [8 s: P# N: X- y"" d4 _. w* F' w% R- D　　二是此卦他是以何爻取的用神？9 v  s+ M2 p( J7 V: M: k& w8 W1 E) \+ K1 L　　三是按癸酉年戊午月乙丑日 湖北某村一男人神秘失踪这个卦语。说明一个问题 他这是先有事发生 了解整个过程 后起的卦。才会有此种情况。. o4 b- o8 x8 ~1 i. X% W5 W"" ?2 {9 K2 [7 A　　他的解释是 从上六起 在兑宫 所以就是口舌引起。牵强得狠。如果他以世爻为用神。那么 与玄武父都不动 构不成关系。* ]% Q4 `9 H% e$ U) h8 P1 M& J0 k5 P1 p) O! r1 a| T* t2 g　　以兄酉金为用 未土来生 也构不成吵架的关系。所以 他这么断 我不认同。& k- M: C! D$ J9 ~- I; v0 x+ c"" p% c　　倒不如动必有因来得直接。% a: V' Z! o/ `- a. d) A  G* b# w+ S$ h' [% j' G0 F9 s　　只看两个动爻 朱雀动 白虎动。朱雀动化出鬼克兄金 由此可知 这是因口舌伤到了兄弟酉金 他临门户 一气之下出了门。+ Q; t4 r* y! c"" g3 m7 \' U3 Q| ]"" a0 E2 ^/  "" K　　此卦因刘文德有一些情况没说清 所以我对有的情况只能从卦中推测。  X) L) w$ K5 G9 U5 z9 p+ h+ C( D* O8 ^'  : ~　　1、从动爻的角度讲 判断出有凶事发生。我认为 他是以世为用神。我是这么看的 以世为用神 父爻为世的克者 所以 断为是他的妻子与他吵架。引发他做出下一步举动"" P| v% b4 k- o7 d8 F* }$ W4 h7 F& N# V% t: Q　　2、父 这个代表妻子的爻临朱雀而动 是口角事。- @2 L7 A/ J8 ]3 `) {. t* q! E3 F0 k( {% p$  　　动化出的官刑克兄酉金。世为阴 所以 顺序从上六开始。上六也是世之财。| K6 }; U- O: w8 A* E5 j! J7 ?' w6 @9 b  q: ~- g6 p　　居兑宫 用神两现 各取所用 它从另一个角度 印证了是口舌而起。' v/ R; ]$ p6 F! E! m8 S- U  T$ p8 S  E2 c+ m　　3、太极转换。未是酒 兄酉也是酒。& v- m3 ?7 K0 }/ k( }/ y/ `0 t: v  C2 Z5 ~+ u# c　　一临白虎 一临玄武。可见 这不是正常的酒。所以定为毒药或毒酒。酉动化退 酉是酒瓶 说明 他没全喝。剩下不少 这样我们就很清楚了。他跟老婆吵架 一气喝了毒药。5 n# R* t+ j0 n4  % M4 Y$ o* O2 K"" L( r& k1 e+ V| E　　4、二五爻均有门户的性质。二是内宅 五是外宅。! D. N! \: {3 g  e4 }; {/ k2 V0 V　　刘文德说：把卦倒过来看 二爻为家 酉为门户 他喝了农药酒以后就离家出了门。我说 不用倒过来 外宅门户动了 临路 所以 他是从家里出去了。从他讲的顺序上说。下一步 应该是到了四爻位。四爻位为蛇 临水 得动爻生 说明是水不少的地方 走到一个曲折的水塘边。' K2 ^$ T! o- @5 Q+ }. L1 W0 `$ }/ k# ?9 \  ~　　刘文德说：泽卦为塘 倒卦的变卦为艮 为东北 所以他出门以后向东北方向的一个大塘走去。因为这里没有山 故艮只作方位论。他从梅花的角度 这么解了一下 我认为 有些牵强。8 U* g' M! q. z5 s2 n: N8 v1 o9 G7 o1 \6 O) l. D　　世爻是卦主。他现在临寅木 居坎宫 这本身就说明了他所在的方面。东北面有水的地方。不用那么费事 硬要把卦随意地乱变来变去的"" ~+ i"" u! @& y7 ^0 G) W% r0 z1 f9 a- D( F　　接着是三爻位了。三爻与四爻位 四之变是午 与三爻位同 是一种接续的方向指引。在这里 刘的论述是：沿着箭头往下看 他的身影已经走到了塘边 这是例卦的二三四爻 是一个互卦的兑卦 兑卦也就是塘。5 ?! B$ N) q$ M: j( ?+ L% f"" u* G& c# r5 V9 X# Z　　二三四是离 二三四变出的是坎 如果按他那么化卦。我看不太懂。: [+ Z! N0 @; B8 f6 ~' D7 {8 {$ t$ V% s; Z; G: L"" x& w　　我直接看爻 四位的水 是到了水边的他 遇见了小鬼。小鬼引着他。让他改变自己 由阳气的寅 变为阴的卯。向死神走进了一步。9 t1  * ]4 R$ F' [) W& e5 `! [2 ?1 f2 j( x# `$ T　　而卯在艮中 是坟地 死人呆的地方。他去了这样的地方- R( d1 t$ f6 i  h+ }1 l# c/ s. s% T0 B7 U6 w　　而午火这个鬼所在的是离火之地 是毒药攻心 动化艮为止 他的生命要停止了。到二爻位的辰土 此土在坎中。土为中央 从另一个角度上 是说他到了水中央。1 @% ~"" d% ]| c. x) @. U9 k/ y' r: B  O8 Z- ~1 ~"" G　　到了水中央 他动了 晃晃当当地 动成了鬼。死了。* o; F! y: ~# C5 T8 s| ~' @9 x8 l| o1 x# M8 i& Z"" h! V2 X) D+ d( s9 o　　四 、巧看外应3 Z% y0 t+ N* O* t% X- V) [; W* H# W4 {6 x　　外应的机理在于把预测时所发现的外界事物作为一种信息 一个兆头 输入到卦中结合而断 有时候可以不看卦而直接就这外应下断语 但更多时候是结合卦来看。因为外应是一种兆象 而兆象本身便是卦象/ S:  2 i$ _# m7 i% L# O|  6 b3  '  + J| l　　外应可以是多个。但这些外应 需要有一个连接性。- ^# s"" C. W' ]$ D* y: @/ z) \: d/ b' M: S( u3 n  E$ y　　外应 说白了 是天人感应的运用。* q$ a6 a# v& M1 w$ W# g8 Q' U  y' C! c0 V8 n| F6 ?; J  v9 k　　（1）卦还没出来 突然出现外应 这个外应可以反映速个这件事的性质 也可以反映事情的开始阶段的状态。0 _1 w0 t8 H* e8 u: L5 a% C2 O; Z4 G8 [　　（2）六个爻全部摇完了 正好在这时候出现了一个外应 这个外应也反映全卦性质。/ V! J3 ~2 c| B! r: y/ {5 _: i; L) o- x7 i# H9 q# ?　　（3）断卦中途出现外应 有可能是应在事的过程中。5 P% L1 E6 i6 O- R/ U| M4 s! `3 `: O| x; y9 O# b　　（4）当写卦至初爻时出现外应 这个外应只反映初爻信息 其它类似。| k' v2 E  u& I' B/ g2 C6 R| B; o% y+ L$ Q　　（5）当我们在一卦中出现几个外应时、要把这几个外应分别对应到与此同步的爻上结合分析"" Q. Q6 @8 u/ m! Z  }3 o5 c' l' C5 w7 o5 ]* m/ A　　如有一次我测算两个篮球队比赛 以甲队为世爻 以乙队为应爻 当摇卦至二爻（世爻）的时候 外面街上经过几辆结婚的喜事车 当摇至五爻（应爻）的时候 恰巧有几只乌鸦从外面叫着飞过 于是即下判断 甲队胜乙队败 卦里面的关系网也不必去分析了。2 d| {3 y/ o# N- G- m. P4 T| ]# D! N! Z& c| ~4 f　　（6）如果一个外应在摇整个内卦时持续存在 那么这个外应反映内卦的事 若持续发生在外卦话 则反映外卦的事。同样道理 持续发生在卦中几个互卦的话 则反映外卦的事。同样道理 持续发生在卦中几个互卦的话 则反映互卦封的信息! J. W; ]3 ~8 q4 s  L; R! t4 X+ z* m3 B　　（7）世爻与应爻是卦中一对至关紧要的座标。当摇至世应两个爻时所出现的外应分别反映世应两爻的事 这种区别对待的政策在预测竞赛 官司 合作 婚姻等二元卦中尤其有意义。| _! {0 y; M& B- S' `& o+ G4 W| J& A| ~* D8 U( N& G# F　　外应与地支、六亲、六神等的结合 建议大家参考梅花三要的应用。比这个更准5 v4 [0 Y  h  D! i7 z' ?4 R  l%  # C$ N5 V! F8 L8 I7 V$ ~2 r0 U　　例一：| M& a) A6 Y# l5 L7 O7 `2 J; j* l9 b1 [$ w　　丁卯年癸丑月丁丑日申酉空 徐先生测生意 夬卦：' k| @$ N| \1 R2 I2 m; Q# b  n6 O$ h) u' _8 l　　　　　　　泽天夬7 ~$ J| r' e% q- ^5 Z% O| B5 Z- z8 d2 l6 F9 J' t　　　　　　　青龙 兄弟未土 ∥/ h5 R7 T0 L' n2 m) A- W4 R) B5 o5 F& H4 ^1 C9 d2 W- K　　　　　　　玄武 子孙酉金 ／ 世9 k- e1 x* k) k& V* P9 c/ Z: m. H0 o4 `  v8 N7 T"" y7 {7 c8 M　　　　　　　白虎 妻财丁亥 ／ 　（有外应）/ Q% r7 {6 y4 H7 w8 f3 x$ i4 P2 e　　　　　　　腾蛇 兄弟辰土 ／: u1 Y9 M; n5 y# z$ M9 Y6 G! u"" N' d! x3 {3 J$ ?* \5 f　　父母乙巳：勾陈 官鬼甲寅 ／ 应! p4 N) @% v"" O: u- G& t0 z( `  z  A8 i# X) {　　　　　　　朱雀 妻财子水 ／- k7 x' \"" C' ?% k6 I2 i( [$ b& ]| T! ?% P　　原断：此卦当摇到第四爻 忽有邮递员送汇款单至 这飞来之财 正好与亥财相对应。亥为猪 于是我叫此人去贩猪肉可以赢利 本来他准备与人合作贩鱼的 听我说了以后 就改变主意去贩肉了 结果赚了大钱。而那位贩鱼的伙计因为路上车子被堵拖延时日鱼都死掉不少 结果赔了本。2 y7 ]3 p; a% u2 }0 e; U  l9 `"" F9 ^# q4 f9 F　　相逢解析：这里 有个先决条件 我们平时在占断时 如果仅凭邮递员送汇款单至 亥为猪就这么断 那么 十有八九 你是蒙对的。1 G) o! `# h0 J; g/  ( v! N' t) q7 H  ]. A　　首先。有汇款 可断为生意得财。' \4 A4 d% ?2 m/ H  h# B+ J"" ~5 N9 K5 c　　但亥水到底是什么财。应该说 鱼他也是水财。不能因为一个亥字 就断为猪了。还要结合其它的象 才能断准: n: h! f8 V1 B% X: S0 J- \& S$ X& l3 ]* b( h| {! [9 r! Z　　其次 此例中 亥水临白虎 显然。老虎样的 鱼不是。猪是这种带毛物。# C& w3 Q) D  O5 k+ u2 i! `8 _* r0 G$ q6 H# D2 J2 d( Y: B　　第三点 在四爻位 与五爻玄武相邻。 一般地 人做鱼生意。不会是在臭水坑中的鱼。 此水居于兑宫 兑为泽。是小水坑类的地方 死水类的。结合玄武、白虎 是不干净的水坑。 而猪是喜欢这样的地方的  通过这样的判断 如果是鱼和猪选一样 才可定为是猪而非鱼。6 I1 X2 g7 ]  C1 S5 i. {5 e' T: }  L- z| I! E　　第四．从卦中的角度讲 此卦的结构不错 但天时并不好。在日月上 是双克亥水。 临财白虎 人在五爻为路。 是做这个路途中的生意钱泄金气 这是赔钱。 结合日月双克 赚不到的。2 S) X8 z) z/ M! ^( m"" t9 a| z| L"" o. ?| M# W　　世临空 说明世主自己心里不托底。应爻官 财生应 还要小心被骗。: N) n. `7 c* ]6 D; Z. r/ ?. w5 d  _1 q/ v　　日月克白虎死猪 世临玄武。而且空 是他要做的这个生意 没经过卫生部门检验 可能是死猪的猪肉。- J( M5 R$ y. h' h1 {6 U0 Y+ M: [1 y- I6 x| V　　如果能得到钱 也是小钱 有欺骗性质的钱。+ c8 ?% M1 K' p"" C# W5 u- T: Y4 V7 O; G% c　　刘文德原断：此卦当摇到第四爻 忽有邮递员送汇款单至 这飞来之财 正好与亥财相对应。亥为猪 于是我叫此人去贩猪肉可以赢利 本来他准备与人合作贩鱼的 听我说了以后 就改变主意去贩肉了 结果赚了大钱。而那位贩鱼的伙计因为路上车子被堵拖延时日鱼都死掉不少 结果赔了本。& ]"" T( _8 X) a1 k; E7 N+ S/ M# O/ K  S7 v/ D6 Z- M( P6 S　　我更相信的是：刘文德断的这个卦的卦主 是做了鱼的生意 赔了本。而做猪的生意 只是他老人家编出来的一个想象中的故事。 如果我编这个故事 我一定会说 他做鱼生意 不听我让他做猪生意的话 赔了本。/ }! K% @& d6 e6 G0 ]: Y+ r8 S* W7 [5 P3 k　　结果 别一个听话的 做猪生意的  赚了钱。这样编 别人就不好看出有假了。9 @4 J- x| E"" w   2 ]% H1 e) d1 b- l# O　　例二：酉年 戍月 壬辰日 刘先生问去南方凭口舌赚钱之事。3 c  O: G) b9 X) U0 `"" x' J: Q: M. U7 B- ^7 j$ L　　　　　　　地火明夷　　　　地山谦' k( n   # x6 u. n' K( i0 R3 E2 \) j  Z  [) i0 L6 c  P6 H- }　　　　　　　白虎 父母酉金 ∥ 　　父母酉金 ∥' ~  D/ F& F. s8 T; n  p9 }9 @4 B' b/ q+ S; X| u5 b5 Z* i' p6 Z　　　　　　　腾蛇 兄弟癸亥 ∥ 　　兄弟癸亥 ∥ 世8 u: E. d0 p: N; A8 q# P% C6 @"" Q  o3 S* ~　　　　　　　勾陈 官鬼丑土 ∥ 世　官鬼丑土 ∥9 Q/ w% t  U/ T1 R1 r5 l2 G; X!  % u　　妻财午火：朱雀 兄弟亥水 ／ 　　父母申金 ／ 　（有外应）+ m' z# p. p! [/ q7 ?- L+ _0 E5 n4 [% m  X　　　　　　　青龙 官鬼丑土 ∥ 　　妻财午火 ∥ 应) b) U8 G. J3 m4 Q3 [# Y- `* U' ]) a4 m　　　　　　　玄武 子孙卯木 ○ 应　官鬼辰土 ∥2 S) w+ [2 `8 Q7 S6 T% p( m- A| }% ]; o2 s　　原断：正摇至第三爻 忽然站在墙上的鹦鹉鸟外型的温度计掉了下来 三爻恰是朱雀临之 朱雀为开口之神。如今这朱雀坠落于地 显然外应不吉 嘴巴饭是吃不成了 更何况卦中飞来克伏 所伏之财又空亡 虽暂有月来半合 但旋即亥月 兄弟值月 财不得出。皆无财利可言。后果在南方跑了十来日空手而归。虽然卦中本有数理之不吉 但这外应鹦鹉临朱雀坠地也是大碰巧了！ 地火明夷已有出行伤人之兆。 测的是求财事 所以 可以应在求财的半途而废止上。 应爻为场所。动化鬼。应入库。动入水库。 没有他施展嘴艺的地方。 财午火出 又入月库  但难出来了。 财不出是无财。' V. Q8 i"" q( c1 a7 n& r3 Z: q- _1 l' f4 D6 ?3 ]7 ?) D+ c  a6 \* q2 d$ o　　世勾陈持 日月双助过旺 说明他嘴里能说的 多是陈词烂调 没有新东西 所以 骗不住人。土持世也主嘴笨。不会说。5 Y0 V/ o9 q; L1 \| n# C# j* X. f4 d) V& D　　看来这是个算卦的 学的是八字 想到南方骗点钱花。9 g' R0 m7 W/ u6 N/ [4 d+ N! P4 m"" W+ l& w9 x6 b' U- V　　外应之所以称之为外应 是因为它具有信息元件的功能 能够称得上外应的 应该具备以下几个条件（这里指动态外应）。! }| m- ^- a* U"" }+ q. v! h9 C# N/ s$ q$ f( v: `0 p　　1、在摇卦的时候出现 无论它是突然的 很快的还是持续的出现 这是指时间上要到位。8 \1 ^/ ~: Q/ D. L0 ]/ h& p3 r8 _$ R　　2、具有一定的象征意义 即具备某种典型性。这是指象的意义上要到位。6 r8 Z7 }! K7 _  Y6 s& x0 W2 ~( g  K"" q- R* c  @2 Q' d　　3、具有一定的力度。外应的力度与事件的程度成正比（如距离远近差别 力度速度差别等等）。.  "" v. e8 i: Z0 l7 U# g* ~"" Y# \5 v: F!  0 `2 \　　五、无中生有; t$ s; w7 I. K! q7 }5 ~: N| i5 B6 x; `  e& R"" o4 o　　六爻卦只有有限的六个爻和地支六亲为六神; z* g* f& \% W"" X& D# l; g1 y. {* _"" J　　卦中还有其它大量的信息存在。9 j8 S| o5 Q. P5 s"" \"" p5 {% O0 b$ {　　“无中生有”基本上有三种表现形式：伏神式；变出式；关系式本文由天机阁 www.tianjige .net 整理  更多内容尽在www.tianjige.net"|http://www.360doc.com/content/15/0215/23/17470473_448876292.shtml|2015-02-16
其他社区|1703641278|kafan|安全&IT资讯|ZHO|2015-03-15 09:01:01|比亚迪欲与特斯拉展开较量 电池产能将增至三倍|据路透社报道 中国汽车制造商比亚迪计划将电池生产规模增至现有的三倍 以此在电动汽车电池供应以及能源储备方面与特斯拉展开较量。比亚迪发言人马修·尤尔杰维奇(Matthew Jurjevich)表示 公司计划 在接下来的三年中 其全球电池产能每年将扩大6千兆瓦时 若需求强劲 公司希望三年后仍按照这样的速度持续增产。这意味着 到2020年初 比亚迪的电池产能有可能从今年年底的10千兆瓦时提升至大约34千兆瓦时。这将使它几乎可与特斯拉投入50亿美元巨资建设的超级电池工厂相比肩。在新兴的电能存储行业中 比亚迪和特斯拉作为两大重要企业正在迅速崛起。储备技术可吸收风电场或太阳电池板的多余电力 并予以存储 留待无法发电的情况时使用 因此被视为整合大量可再生能源的关键因素。比亚迪美国分部的尤尔杰维奇在采访中表示 “我们已经证明 若市场需求强劲 比亚迪有能力每年增产6千兆瓦时。”电能存储行业吸引了特斯拉、比亚迪以及众多初创公司乃至一些大型电池制造商。市场研究机构GTM Research预计 单独美国市场而言 到2019年 这一行业的规模预计将从2014年的1.28亿美元攀升至15亿美元。比亚迪的生产主要集中在中国 但今年还将在巴西开办一家规模不小的新厂。尤尔杰维奇透露 该厂将为明年的产出做出巨大贡献。由于电池需求不断在增加 比亚迪也将扩大公司在美国的生产规模。据市场研究机构Lux Research去年发布的数据显示 比亚迪是混合动力汽车和插电式电动汽车的第六大电池制造商。为特斯拉制造电池和电池组的松下则位列首位。特斯拉当前虽不生产电池 但在2016年 该公司将在内华达州启动电池生产 直至2020年 其产能将达到35千兆瓦时。2013年 比亚迪在加州南部开办了两家制造工厂 生产用于公共交通的电动巴士以及电池。比亚迪在2003年开始展开汽车业务 这在当时令业内颇为震惊。此后 该公司已成为中国最成功的汽车制造商之一。但在国外 比亚迪主要销售巴士而非汽车。在美国 比亚迪计划今年部署70兆瓦时的项目 另外还有130兆瓦时的部署计划仍在筹备中。在北美 已有40兆瓦时的项目部署到位 其客户包括雪佛龙(Chevron)和杜克能源(Duke Energy)。(陈思) 随机推荐 今早更新307要求重起！  请问浪滔天的汉化哪里有下？  高手们请帮忙！！！ka60激活问题v7&period;o&period;o  关于Returnil Virtual System和Returnil 虚拟备份7版本争执  关于局域网内ARP攻击源的问题  avast主页的那个有图案数字的金属圆球是神马？  Immunet 卡饭admucher ipv6windows 2003 server 杀毒ess6&period;0&period;316更新慢indesign cc 64bit baidur studio7&period;6注册码parite 病毒eset nod32 server2003mdk3 下载接收的qq文档不显示图片|http://bbs.kafan.cn/forum.php?mod=viewthread&tid=1816113&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline|2015-03-15
기타|1703730943|ngzb|新闻互动|ZHO|2015-03-15 10:51:01|说好的“变形金刚”、“梦幻海洋”、“神秘森林”呢?南宁一气球展被投诉与广告不符|"马上注册 结交更多好友 享用更多功能 让你轻松玩转南宁您需要 登录 才可以下载或查看 没有帐号？立即注册  x说好的“变形金刚”、“梦幻海洋”、“神秘森林”不见踪影南宁一气球展被投诉与广告不符0 X# [+ C# v5 f; q　　南国早报网―南国早报南宁讯 （记者经小飞）3月14日 很多家长通过商家网络广告慕名带孩子到南宁市凤岭儿童公园看气球展 发现商家广告中的“变形金刚”、“梦幻海洋”、“神秘森林”等造型压根没有 而只有一些简单的气球造型。不少市民带孩子进去转几分钟就出来了 并大呼后悔来看。+ ?8 K5 ~"" u% Z9 U( f3 N: V% m"" u"" d2 J　　近日 一则“南宁市凤岭儿童公园周末有气球展”的广告迅速在微信朋友圈传开 原来 商家承诺 只要到售票处出示转发此广告的记录 即可享受半价20元。广告的图片中 有“变形金刚”、“梦幻海洋”、“神秘森林”等大型气球造型。市民翟女士收到了朋友分享的这一信息 便于3月14日带孩子前往观展 不料现场只有十多个简单的气球造型 整个展厅“就像一个大仓库” 几分钟就看完了。她一出来就在网上发帖 大呼失望。5 ?0 l| d' S6 A. a' Q% Y+ M: P1 q2 H+ q4 P6 Y　　接到反映后 记者于3月14日下午来到凤岭儿童公园举办气球展的梦幻城堡。现场有上百人排队买票 非常热闹 不少排队的家长都说是被朋友圈转发的广告吸引来的。( D( Z3 R$ o! g  [0 r( O| m4 q1 W* ^& h$ L% ^　　记者花20元钱买了一张门票入内 只见气球展设在一个约500平方米的展馆内 场内共有13个气球造型 有彩虹、海绵宝宝、机器人等 造型相对简单 规模也小 广告中的“变形金刚”、“梦幻海洋”、“神秘森林”等大型造型不见踪影。展馆光线很暗 走一圈 几分钟就参观完了。有的市民还是从西乡塘专程带孩子赶过来看展览的。记者随机询问了10名进去参观的家长 他们均表示 气球展的实际情况和广告相差太远 这20元门票钱冤了。0 T"" g| K1 O2 F| J2 r% R1 \: h. ?- L　　为何现场的气球造型跟商家广告宣称的不一致？售票的有关工作人员解释称 广告上的图片是在其他地方展出时做的 因展览场地不同 造型自然不一样。/ ]0 ~6 Z: x; n7 K9 V% E  ?"" I4 ^. m　　凤岭儿童公园服务科的有关负责人表示 为丰富儿童公园的活动 在气球展览公司的建议下 该公园联合对方举办了气球展。由于在做广告时 展馆内的气球造型还没做好 因此用了以前做的一些造型 加之城堡内展出的面积不很大 考虑到游客参观和孩子拍照等问题 故造型和规模均有限制。而且气球的造型要根据不同的展出场地来打造 他们在广告时也就此作了说明。该负责人也说 因气球造型都是纯手工活 做起来很不容易 因此不能简单地用“值不值”来评价。对于观众提出的意见 公园深表歉意 也会进一步跟气球展主办方沟通 争取再多制作一些气球造型。) R7 c. ~3 j* E; u' m2 `) L7 G1 k3 V( Q! @0 w7 S. T　　（读者某女士 稿酬50元）& @/ k8 C- ?% R6 v8 u5 o* @3 l$ E$ i) ]'  - H3 l4 d  a2 G8 Z南宁| 气球展| 被投诉| 与广告不符"|http://www.ngzb.com.cn/forum.php?mod=viewthread&tid=922081&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline|2015-03-15
기타|1705050629|ngzb|新闻互动|ZHO|2015-03-16 10:49:01|3・15携手共治 畅享消费：央视3・15晚会曝光多家企业|"马上注册 结交更多好友 享用更多功能 让你轻松玩转南宁您需要 登录 才可以下载或查看 没有帐号？立即注册  x央视3・15晚会曝光多家企业8 v2 q* O; A7 }5 F| V登录/注册后可看大图17.jpg (25.25 KB| 下载次数: 0)下载附件 保存到相册25 分钟前 上传</ignore_js_op>内幕人士爆料。: R- ?. j| l+ t! j　　东风日产、上海大众、奔驰4S店：$ q* q  e& N# d  [$ h; A8 x% E　　小病大修 牟取暴利+ x. l5 e! ~* w' J% y$ s; ^. a% R1 g8 e5 ]5 x1 u( V$ ^　　记者调查4S店发现：东风日产、上海大众、奔驰4S店会故意虚报和夸大车辆故障 从中牟取暴利。一辆简单故障的汽车（点火线圈插头松动 重启系统即修复） 在这些4S店 却要你更改火花塞等各种大修 其中奔驰维修费报价近万元。/ Z) m; B;  8 j# Q! E0 B$ w8 S' G( E! Y　　央视3・15晚会节目组接到了大量消费者投诉 纷纷反映一些4S店在车辆维修和保养的时候 存在许多猫腻。一位多年从事汽车维修的内幕人士 也向节目组举报 一些汽车4S店会故意虚报和夸大车辆出现的故障 欺骗消费者 从中牟取暴利。8 q9 T; w! x/ b. u$ O5 d5 I6 t6 h  J- D: a5 H; n& J& g% b　　内幕人士告诉记者 一些4S店常用手法是“小病大修 没病大修 能换的不给你修 能修好的也要求给你换”。* r5 F% ?7 m7 @0 {(  7 j| v6 n* ]/ H4 M2 b: I3 l) e　　真的像内幕人士说的这样吗？记者决定对4S店的售后服务进行调查体验。) `( I6 O* ~- }/ P; v+ a; \) O* R8 ^. d1 c　　这次体验调查 记者设置相同的简单故障 在北京、天津、河北、河南、安徽、上海、浙江等七个省份 先后22次对东风日产、上海大众以及奔驰的4S店售后维修进行体验调查 遭遇小病大修的次数高达16次 比例占到73%。) V( K# U6 e& A' u* p( i4 C+ F+ E4 \5 r| p"" f' W　　路虎成恐怖的“拦路虎”% `: ^- D( q3 B3 a3 R$ ~$ M* h7 M# F0 _6 w5 d+ t　　说起路虎揽胜极光车 消费者用最多的词是“恐怖”。要么走在路上不动了 要么倒档失灵 全国类似案例不计其数 虽然这被诊断为变速箱故障 但部分车主说换了两次变速箱仍故障频发。路虎中国公司甚至将变速箱故障原因直接推到用户身上 嫌车主开车太着急。3  ( r2 }) N8 X) ^* Z5 `6 V8 Z% N$ @5 X( r　　宁波杨先生这辆路虎极光车在倒车的时候 故障频发。“就是R挡（倒挡）一直闪烁 然后我踩油门 看到没有我就是加到红色了 车子都不会动 一点都不会动。”2 p5 _1 m! p5 I) j3 K5 R% s! B; l! D　　在宁波路虎4S店里 杨先生遇到了因同样问题来维修的车主冯先生。2 a& p1 S' @7 F. h* m( i0 m' T9 D/ r% W! _8 f　　冯先生的路虎极光车刚开了两个多月 这已经是他第四次去4S店了。“一挂倒挡车子往前冲 不走了 怎么挂挡也没有用。”- P/ U; U2 k8 I  d+ u9 ]/ }* J$ ]& E1 j9 N| m4 m　　记者了解到 路虎极光是路虎旗下一款进口豪华城市SUV 2014款和2015款配备了9速自动变速箱。然而 出现严重故障的 正是这款路虎极光引以自傲的9速变速箱。: U% @! P# D+ R# ]+ K/ T3 a# _; j6  (  "" Q- z; i1 H　　软件升级是路虎公司针对变速箱故障给出的技术解决方案 不过 路虎4S店很快发现 这个方案根本无法解决频发的变速箱故障。/ h( X; Q( V6 n0 C$ f. z/ B& D"" I' G+ ^4  ! R. K9 [　　北京刘先生的这辆2014款路虎极光车 在软件升级后还是多次出现故障 最后不得不更换变速箱。; c4 _0 Q$ k- R4 ~$ }1 H0 y$ j3 h5 K( A- ?$ M- O; c"" B' c　　虽然给出了方案 但对于变速箱故障 路虎中国始终不愿承认。在路虎中国的官方网站上 记者始终看不到任何关于路虎极光变速箱故障的说明或者公告。/ l% U; S1 Y$ c# M# o; `: u$ @3 P% M; ~"" L. h　　面对越来越多车主的质疑 路虎中国公司却将变速箱故障的原因 直接推到了用户身上。捷豹路虎汽车贸易（上海）有限公司工作人员称 是国内车主开车太急了。  l0 \. Z) H* ^4 U7 H& U"" ]"" P+ H/ a8 M) G. X　　车主们想知道 车辆一旦过了保修期 谁来承担变速箱故障带来的高额维修费？更让车主们担心的是 因变速箱引发严重的交通事故 谁来为他们的生命安全负责？; k/ H6 ]| [$ S4 j) P/ C5 e| }' e* K"" w  F　　山东不法厂商调和有毒汽油0 c8 h3 Q9 k4 N  e8 Q7  8 y% z4 P9 _　　加油后车子还没劲、抛锚？真相：在山东省东营市、滨州市许多不法厂商调和各种石化原料 年产量达五六十万吨 获取暴利！而且！这种调和汽油竟然还符合国家标准 加油站默许直接加到了咱消费者的车里 调和汽油含甲缩醛 易造成汽车线路漏油 还会挥发有害气体 污染环境 影响健康……| S/ W| o- @' k2 m) d8 s( @' u1 r! ?7 F2 P　　最近全国各地的许多车主反映 他们的汽车加油后会出现没劲甚至趴窝的现象 怀疑汽车出了问题。一位业内人士向记者曝出了其中的秘密 问题就出在了汽油上。一些不法厂商通过调和各种石化原料 大量制作出所谓的调和汽油 获取暴利 而各项指标检测还完全符合国家标准 在加油站更是一路绿灯 直接加到了咱消费者的车里。"" u# i* L8 i1 C# x:  . p: T7 K6  | ?/ G- ]4 u4 p　　记者连续走访了东营、滨州等地的多家生产调和汽油的工厂后发现 这些企业大部分都用石脑油、抗爆剂以及其他一些化工原料做简单混合后生产调和汽油 价格比正规汽油便宜很多 销量可观 并且这些企业负责人都信誓旦旦地声称 他们生产的调和汽油都能符合汽油国家标准。因为现行的汽油国家标准中规定 只要通过辛烷值、硫含量、苯含量等十几项检测标准就判定为合格的汽油。至于汽油里具体含有什么样的成分 并不在标准的检测范围之内 这就为调和汽油生产厂家带来了可乘之机。& I+ M) ^! ]6 O: L! s( P! f; c* e5 S1 V% p7 @- J"" D* F% i1  　　记者调查发现 在山东大大小小的调和油厂就有200多家。. M7 p0 x/ i& n& B5 d* J3 Q' Q  U# A+ n/ ?　　甚至还有人开起了培训学校。淄博圣通化工研究所虽然挂着研究所的牌子 但主要业务却是调和汽油的培训 三年来已经办了90多期培训班 为全国各地培训了800多名技术人员。! i) t; _$ y8 U0 X: Q  m9 Q& m* K2 v( ]0 H4 M"" C　　电讯企业成诈骗电话幕后推手% \! V) z- Z& r- a1 p6 ]0 ~* N0 i: {. v3 L( e% O　　骚扰电话 有时一天要接好几个甚至十几个 对方有时候还冒充警方、银行等诈骗 谁是它幕后的推手？你肯定不敢相信 中国移动、中国铁通在为骚扰电话提供各种支持 甚至给“10086、110”之类的诈骗电话一路开绿灯 及时发现诈骗电话显示虚假主叫号码 仍然允许透传。; C# }& q1 i0 ]9 x  H$ T) Y8 W% q4 w. h　　群呼电话、显示虚假电话号码 不仅为骚扰电话大开方便之门 更是被一些不法分子所利用。大量公开报道显示 不少骗子正是利用了群呼、透传等技术 将主叫号码显示成银行、公安局、法院等单位的电话号码实施诈骗 诈骗金额少则几百上千 多则上百万。7 f/ ]- j8 e| B% o2 {# m) F0 Z+ x; \. _7 I/ R5 B9 ?　　在运营商的默许和技术公司的大力支持下 呼叫中心将越来越多的电话拨给了用户 而我们也只能一次又一次地被骚扰 一次又一次地被动应付。/ `4 U* ~4 j$ Q2 a- }2 R# S2 e2 }! t( h7 R- R6  8 l　　手机实名制形同虚设：随意买到电话卡; F0 y. q"" m8 S7 i  H| @8 f: S| X: v6 q% ~| _　　记者调查发现 联通公司员工为完成开卡任务 偷偷利用消费者留下的身份信息 再次重复激活开卡（一身份证可开五张卡） 完成开卡任务 余下手机卡20元/张卖给卡贩子 卡贩子卖给诈骗犯。你名下有没有手机僵尸号？小心有天警察找上门。6 ^"" `% @8 j: k% ^$ J7 I0 `# V| L/ k6 N5  ( S' I　　银行存惊天漏洞：你正沦为洗钱帮凶"" [. \5 t- z4 z' X"" J& {1 P* y0 E4 R+ n　　诈骗犯到底咋洗钱？他们从网上购买一套真的身份证+银行卡+手机电话卡=成功用此转移财产。那么问题又来了 这些银行卡哪来的？记者深入调查发现惊人内幕：网上买一张别人丢失的身份证 拿去四大银行 其中工商银行、中国银行、农业银行可轻松办理银行卡。' U5 B- X"" l  E1 h0 z6 y! H  `$ e' Y8 {; o( q/ p: M| y　　记者发现在一些QQ群里 有人在公开兜售身份证和银行卡。在一位卖家的QQ空间里 几百张身份证被拍照上传供买家任意挑选。每张价格200元左右。这名卖家告诉记者 他每年能够卖出四五千张身份证 其中大部分被用来办理银行卡。不仅身份证公开买卖 甚至连同用身份证开户的银行卡也可以成套出售。在网上像这样公开买卖身份证和银行卡的QQ群 可以轻松地找到几十个。* e"" r. k; J$ B+ y  s3 k| [' J8 q% z  C: s+ Z) W' t4 y% {5 O　　随后 通过一名卖家记者购买了 工商银行、农业银行、建设银行和中国银行四套银行卡。+ p1 I7 q/ R3 y( e' F: ]: ~! `% H| w+ }  G| ~　　这些银行卡 除了开户人的身份证以外 还包括网银U盾和绑定的联通手机卡 经过测试这些银行卡的网银、转账、支付等功能一应俱全。5 o0 Q8 u9 g4 f  K3 ~% a! J! j6 p　　那么这些功能齐全的银行卡究竟是怎么办出来的？根据国务院颁布的《个人存款账户实名制规定》 个人在金融机构开立个人存款账户时 应当出示本人身份证件 使用实名。- L6 U: @& e$ J# D+ A1 `5 z9 j4 Y) A( k3 V0 W7 b& M5 p) u4 b　　用一张买来的身份证 在北京工商银行西四环支行 工作人员没有任何疑问 记者就顺利地办出了银行卡。+ Z& r% Z2 G9 X7 y) S) f* n& v) B' y  r# c' e　　在中国银行和农业银行虽然工作人员也发现身份证上照片与记者明显不符 但记者还是顺利地办出了银行卡。& A0 W( e3 O( ?3 Q+ k; i1 W: I4 m"" H　　仅凭一张从网上购买的身份证 记者就轻松地办理了三张功能齐全的银行卡。( x. b$ A' }0 \2 w4 \4 m4 e| }$ }/ v+ q6 V/ G　　正是利用银行这个漏洞 网上一些人专门帮助骗子干起了洗钱的勾当。一次洗钱的过程会涉及到几张甚至几十张这样的银行卡 这也给警方追缴受害人钱款带来极大的困难。! o: E"" }  [' l7  1 \9 k6 T! I8 l1 Y$ N| v5 D!  + x　　深圳保安分局网警雷耿告诉我们：“他们买的这些银行卡 如果追查的话 基本也就是追查到开卡人这一级 用卡人这一级就很难追查。”9 `3 e- t+ [* d' T5 D& b% D# G5 K' k3 l& f0 j. g; O#  　　就这样 这些在网上随意买卖的身份证和银行卡 成为一些不法分子大肆骗钱的有利工具。1 E7 {1 A: A| P4 G. N: H-  ; v6 t"" v7 ~; {; A3 H) q$ s( y　　谁来管管来路不明的保健品？6 t/ O3 F3 B( J1 \| i3 F! v4 r; q2 i+ ]6 T3 I1 k6 ?$ s( c　　72岁的王大妈 平时省吃俭用 为了健康 偏爱购买各种保健品 在她家里大大小小13个纸箱子里装满了这几年买的部分药品 总共有30多个品种 投资近40万元。但记者仔细看了看这些所谓的药 大都没有任何批准文号 来路不明。王大妈怎么都不相信 保健品并没有给她带来健康 留下的除了一身的病痛就是沉重的外债。7 C7 i; L; R3 l& }; j9 `( ?8 ~3 V- a$ w. l　　记者在采访中一再提醒王大妈 不要再上当受骗。可是 大妈已经深陷骗局 不能自拔了。当记者第二次去采访王大妈时 她又买了一个艾灸治疗仪。可恨的骗子榨干了老人的养老钱 留给大妈的只有虚幻的健康。其实 这些不法商家是怎么忽悠老人的？总结惯常的骗术 有四招：4 O2 W5 @) ~: l. }8 ^| X. {"" O/ b- s& K0 N% z# Q5 b2 h　　第一招 洗脑营销。打着免费健康讲座的旗号 向老年人灌输歪曲的健康理念 虚构夸大他们的病情 诱惑老人买保健品和治疗仪器。3 U9 v$ }! V# u; {) E! Y4 W3 w4 m* e2 r% B2 G! x　　第二招 亲情营销。营销人员一见面就喊爸爸妈妈、爷爷奶奶 哄着老人高兴 其实看中的就是老人兜里的钱 让他们最后买了保健品。"" a* U9 ?$ O1 p6 z2 q8 {* p$ w& E  q0 n"" Z9 l8 U5 v　　第三招 体验营销。拉着老人体验各种医疗器械 吹嘘疗效 忽悠老年人花钱。  m3 W' t; n& u1 g# V2 o"" }7 S7 Q9 E! l5 ]| U　　第四招 免费体检。打着免费体检的幌子 在体检报告上做手脚 吓唬老人赶紧掏钱治病。( a4 k$ r8 n( a2 }$ C2 D/ G2 j( N9 p0 B- r6 z　　央视3・15晚会截选报道6  2 I& O+ r7 }6 s3 u# \% a& M0  + F2 j; ^1 k+ w( p/ U1 p2  + d( {% U' S| W2015| 央视3・15晚会| 曝光| 多家企业"|http://www.ngzb.com.cn/forum.php?mod=viewthread&tid=922226&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline|2015-03-16
其他社区|1729423167|360wenda|已解决|ZHO|2015-03-31 12:01:01|朗逸13款1.6l自动豪华和14款1.6l自动运动哪个好|"个人建议你选择14的这款 相对车型较新 技术更加成熟 其实你看中13那款无非是内部配置而已 如果仅仅因为这个 建议你还是买14这款 毕竟降价处理的东西总有在年份上的缺失送给回答者一份礼物送香吻 赠言：好帅的回答 楼主送上香吻一枚 以表诚挚谢意！ 00x用微信扫描二维码分享至好友和朋友圈分享到：检举 -->答答好搜问答团队最勤劳最可爱的答答15分钟前下面是答答童鞋给您的小建议 您看靠谱吗？初来乍到 弄错了您不要生气哦(*^__^*)答答小贴士相关问题13款上海大众朗逸1.6L自动舒适版和广汽本田凌派1.8L豪华版哪...12014.03.2113款迈锐宝2.0自动豪华、新朗逸1.6自动舒适哪个费油呢。上下...2013.11.15k315款1.6l自动dlx和朗逸13款1.6l自动舒适版哪个好2014.11.24英朗GT1.6L自动舒适版和新朗逸 1.6L 自动豪华版哪个好呢|求推...122013.09.10朗逸13款自动豪华和改款的区别2014.11.22查看更多关于的问题 >>"|http://wenda.haosou.com/q/1427769875725878|2015-03-31
其他媒体|1729912520|tieba_baidu|Keyword_笔记本吧|ZHO|2015-03-31 17:22:02|《盗梦英雄》3月庆公测 抽大奖 送豪礼！|这个活动很给力 小伙伴们不要错过哦！来自: 盗梦英雄官方  -盗梦英雄吧时间：2015.03.19 - 2015.03.31状态： 活动进行中奖品： 京东礼品卡100元、《盗梦英雄》限量定制抱枕、《盗梦英雄》限量定制... 动态： kapdxi813619获得了《盗梦...  -7小时前  xt523188获得了《盗梦英雄...  -7小时前  sleepdian81获得了《盗梦英...  -7小时前  kuatoe231获得了《盗梦英雄...  -7小时前  mataoohye88116获得了京东...  -7小时前  *********获得了《盗梦英雄...  -7小时前  shoujjjio获得了京东礼品卡...  -7小时前  sc4Me8688q3w获得了《盗梦...  -03-25  zhou081获得了《盗梦英雄》...  -03-25  3n1ri23n74bp9t获得了《盗...  -03-25  jinboyiyi获得了《盗梦英雄...  -03-25  apm1861获得了《盗梦英雄》...  -03-25  kemeng30118获得了京东礼品...  -03-22  SEC研获得了《盗梦英雄》限...  -03-21  空白格LV1获得了《盗梦英雄...  -03-21  一枝花大姐获得了《盗梦英...  -03-21  净石123获得了《盗梦英雄》...  -03-21  九年义务631获得了《盗梦英...  -03-21  酒徒_ze获得了《盗梦英雄》...  -03-20  花妖娜娜228获得了《盗梦英...  -03-20  时尚假发专门店获得了《盗...  -03-20  wnk3i1mdxo7m5q获得了《盗...  -03-20  tutu486966获得了《盗梦英...  -03-20  月冷枫清谈获得了《盗梦英...  -03-20  他就是先帝啊获得了《盗梦...  -03-20  *********获得了《盗梦英雄...  -03-20  邓家柒少获得了《盗梦英雄...  -03-20  袁书华2008获得了《盗梦英...  -03-20  钟凝2获得了《盗梦英雄》豪...  -03-20  一片叶2046获得了《盗梦英...  -03-20  淡淡烟草味0409获得了《盗...  -03-20  zhuqin*******获得了《盗梦...  -03-20  蝶舞嫣蕾获得了《盗梦英雄...  -03-20  *********获得了《盗梦英雄...  -03-20  遗忘浪子520获得了《盗梦英...  -03-20  麦兜来来来获得了《盗梦英...  -03-20  冰毒之ICE获得了《盗梦英雄...  -03-20  坚强的小志获得了《盗梦英...  -03-20  tuyuan********获得了《盗...  -03-20  北交大迎风而立获得了《盗...  -03-20  tulin_2获得了《盗梦英雄》...  -03-20  会会飞飞飞飞飞获得了《盗...  -03-20  郭建忠888188获得了《盗梦...  -03-20  阿拉420获得了《盗梦英雄》...  -03-20  大肥超2013获得了《盗梦英...  -03-20  蒸发眼泪1013获得了《盗梦...  -03-20  tuwen1010获得了《盗梦英雄...  -03-20  苏是我媳妇儿获得了《盗梦...  -03-20  漫无边际1970获得了《盗梦...  -03-20  v任逍遥0获得了《盗梦英雄...  -03-20    立即参加 15.5万人已抽奖|http://tieba.baidu.com/p/3670673113|2015-03-31
各大媒体|1744217673|news_baidu_search|search_现代汽车|ZHO|2015-04-09 16:26:02|起亚k3和朗动哪个好 北京现代朗动2015款 朗动全系低价促销|"来源:汽车中国 作者:匿名 发布时间:2015-04-09 [查看评论]<\/a> 关键字:低价 促销 北京现代 哪个 1.6L 朗动的内饰有着明显的家族特征|颜色搭配也采用了..."|http://new.carschina.com/jinkouxinche/201504091270624.html|2015-04-09
汽车社区|1745420026|sina|国内 > 最新消息|ZHO|2015-04-10 10:21:01|深度：枭龙战机如何参与也门空袭 做对地攻击机|　　　近日 巴基斯坦枭龙Block2战机的总装线曝光 巴基斯坦方面声称“枭龙”/超级雷电JF-17 Block2战机有多处改进 如航程有所增加、改进雷达、增加探测距离、增加超视距攻击能力、可携挂各种确制导武器 并加装了空中受油管。另外巴方称年产量将从16架逐步增加到25架。　　新浪军事编者：为了更好的为读者呈现多样军事内容 满足读者不同阅读需求 共同探讨国内国际战略动态 新浪军事独家推出《深度军情》版块 深度解读军事新闻背后的隐藏态势 立体呈现中国面临的复杂军事战略环境 欢迎关注。　　近日有消息说巴基斯坦空军将派出JF-17战斗机参加以沙特为首的多国部队空袭也门什叶派武装 这将是JF-17的首次实战。　　由于也门什叶派武装缺少空中作战力量 虽然有消息说他们缴获了数架政府军的米格-29战斗机 但是没有完善的指挥引导、后勤保障系统支持 这些战斗机能够发挥的作用也不大 所以JF-17更多则作为对地攻击机来做用。　　众所周知 巴基斯坦空军由于规模有限 一直要求自己的作战飞机具备对空和对地双重作用能力 这样能够以较小数量的作战飞机执行更多的作战任务 在印巴战争之中 巴空军曾经用F-86战斗机突袭印度装甲部队 阻止了对方前进 协助地面部队有效的巩固了防线。所以巴基斯坦也要求JF-17是一种能够执行空战、对地精确攻击、反舰任务的多用途作战飞机。国产WMD-7光电瞄准吊舱　　对地攻击 尤其是打击地面小型目标首先解决的就是对地探测问题 在过去在昼夜复杂条件下探测地面小型目标是一个难题 比较典型的系统就是美国的蓝盾系统 它由全天候导航吊舱和光电瞄准吊舱组成 此次参加空袭的沙特空军F-15S战斗轰炸机就配备有这样的系统 不过美国出售给沙特的简化型系统 全天候导航吊舱取掉了地形跟踪雷达 后者则取消了发射AGM-65小牛导弹的能力。机载APG-70的对地模式也有所简化。　　JF-17配备的KLJ-7脉冲多普勒火控雷达 它拥有较多的对地工作模式 包括多普勒波束锐化(DBS)、合成孔径成像(SAR)等高精度对地攻击模式 其中后者是利用信号/数据处理系统“合成”一个较大的天线孔径 以提高机载雷达的对地分辨能力 它解决了机载火控雷达探测地面小型目标的问题 还具备地面移动目标指示能力(GMIT) 这样战斗呆账就可以在昼夜全天候条件下探测地面小型目标 提高战斗机的对地攻击能力 所以我们看到新世纪机载火控雷达一个升级项目就是配备SAR模式。　　SAR模式还为另外一种武器的使用提供了便利 那就是JDAM SAR模式探测到目标之后 飞机可以把目标坐标传递给JDAM 然后投掷炸弹对其进行攻击 JF-17配备了我国第一套激光惯导系统 并且整合有卫星导航接收机 可以为飞机和精确制导武器提供高精度目标坐标 JDAM方面巴基斯坦已经从我国引进了FT-2型INS/GPS制导炸弹 并且实现了国产化 这样就可以经济、快速为巴基斯坦空军提供了一种精确打击手段。JF-17挂载WMD-7想像图　　JF-17飞机员可以利用机载火控雷达的SAR模式探测地面目标 利用机载导航系统为其进行目标数据装订和初始对准 然后投掷炸弹攻击目标 不过目前我国北斗二期工程还没有覆盖中东地区 FT-2在也门投放只能使用GPS信号 尽管美国对于此次空袭行动持支持态度 但是FT-2肯定无法使用高精度的P码GPS误 只能使用较低精度的C/A码GPS信号 这样它的投放精度会受到影响 不过依然可以得到从普通炸弹高许多的投放精度。　　对于他国空军使用JDAM这样的武器来说 一个受制于美国的GPS信号 投放精度也不如激光制导炸弹 还有就是JDAM目前攻击移动目标比较困难 所以许多国家空军在战斗机配备光电吊舱来弥补这个不足 JF-17配备有我国WMD-7光电瞄准吊舱 它安装有前视红外探测系统、CCD摄像机、激光测距/目标照射系统等 WMD-7可以在昼夜全天候条件下为战斗机提供地面/海面目标搜索、识别和跟踪 并且对目标进行标定和照射 为激光制导炸弹提供制导 并且还可以提高普通炸弹的投放精度 WMD-7还具备一定的空空目标跟踪和辅助导航功能。它对于地面小型目标如坦克 可以提供20公里左右的探测距离 配合激光制导炸弹 JF-17具备了在昼夜全天候条件下打击地面低速移动目标的能力。　　巴基斯坦方面声称“枭龙”/超级雷电JF-17 Block2战机有多处改进 如航程有所增加、改进雷达、增加探测距离、增加超视距攻击能力、可携挂各种确制导武器 并加装了空中受油管。另外巴方称年产量将从16架逐步增加到25架。　　当然激光制导炸弹也有自己的不足之处 就是受天气影响较大 尤其是也门这样沙漠面积较大的国家 沙尘、烟雾对于激光尤其有影响 而JDAM的优点就是受天气影响较小 所以在伊拉克作战的美军战斗机会混合挂载这两种武器 甚至还出现了混合JDAM、激光制导系统的激光-JDAM复合制导武器。　　对于JF-17来说 由于空中威胁较小 它可以将主要载荷、挂架用于空地武器 如在机翼和机腹各挂载一个副油箱 翼下挂载2枚FT-2型500公斤级精确制导炸弹 翼尖挂2枚PL-5E-2空空导弹 以应付可能出现的威胁 在这种情况下 其作战半径可能达到700公里 足够支持从沙特南部机场起飞 打击也门首都萨那 如果想混合挂载FT-2和激光制导炸弹 这个时候飞机的挂载可能就要变成机腹挂WDM-7 机翼下各挂一枚FT-2和500公斤级激光制导炸弹 作战半径就要受到影响 可能需要从吉赞这样靠近沙也边境的机场起飞 吉赞机场距离也门首都萨那的直线空中距离在250公里左右。　　因此对于巴基斯坦空军来说 今后会把现役的JF-17加装空中加油系统 以提高他们的航程和作战半径。(作者署名：鼎盛军事 小飞猪)　　《简氏防务周刊》称：Block2型JF-17战机安装的是KLJ-7型机载脉冲多普勒火控雷达 图片拍摄于2月19日 这是巴基斯坦航空工业公司生产线上的几架战斗机之一。目前正在研制的block3型战机 将会安装新型的有源相控阵雷达（AESA）。　　本栏目所有文章目的在于传递更多信息 并不代表本网赞同其观点和对其真实性负责。凡本网注明版权所有的作品 版权均属于新浪网 凡署名作者的 版权则属原作者或出版人所有 未经本网或作者授权不得转载、摘编或利用其它方式使用上述作品。 　　新浪军事：最多军迷首选的军事门户！|http://mil.news.sina.com.cn/2015-04-09/1643827314.html|2015-04-10
汽车社区|1859411110|autohome_cn|智跑论坛|ZHO|2015-06-18 00:32:01|老爸购车。车友戳进来|2015-6-17 23:24:05   来自 汽车之家Android版    老爸购车。车友戳进来        话说老爸看汽车之家已经好几年了 他很喜欢车 但是身上没米所以买车的想法放了好久。老爸是个工薪阶层 没多少存款 首付要靠亲戚借来 之后是银行贷款月供大概要在2500左右可以接受。――――――――――――――――――――――――――――――――分割线――――――――――――――  ――――今年爸不知道怎么犯车瘾 非说要买辆开。于是上汽车之家看车来了 一开始的时候是说要订福特福克斯但是因为空间和油耗放弃了 然后是各种看起亚k3 本田凌派。后来感觉家里人多又经常下乡所以看上了suv 在4s看了本田xrv和缤智。可万恶的4s店一分不少还有必须订一万的装修费并且要等一个月提车果断pass。无意间看到新款15智跑gls本地降价2万后16.88万 瞬间的好感啊 立即打电话去了4s导购说在做活动到现场还有东西现车大大滴有。因为舅舅就是智跑高配的还特地花了两万换轮胎 做过他的车感觉很不错在路上开的挺稳的。给爸看了下 智跑的配置爸是完全看好 估计如果米够的话直接上智跑了。  本人初二狗 爸快40了。他的第一辆车我觉得必须帮他选到不后悔 智跑正在考虑 看了很多的车感觉智跑性价比没得说。最后求车友门给个祝福吧。      用户名   操作   操作时间   查看全部|http://club.autohome.com.cn/bbs/thread-c-2137-42511787-1.html|2015-06-18
其他社区|1860230395|yam|即時 > 宅趣|ZHO|2015-06-18 13:21:01|北韓《高麗航空》飛機餐　時隔三年餐點有變化嗎？|圖片來自：instagram.com/jonoh高麗航空在眾多航空公司中一直是獨樹一格的存在 因為國情的關係高麗航空在制服上略顯保守 雖然之前已推出新的航空制服 但整體感還是與其他國有所差異(不過這也成為北韓的特色之一)。當時除了介紹高麗航空的紅藍制服外 還有順道分享讓遊客稱奇的飛機餐 他們家的飛機餐一樣秉持獨樹一格的特色(誤) 以至今日還是有遊客拿出來討論。  高麗航空的深藍色典雅制服 圖片來自：facebook.com/dprk360原汁原味的內容在這裡 原本大紅的空服換成沉穩的深藍 偏高領... 【文章內容不代表蕃薯藤立場 想看更多歡迎到>>>卡卡洛普－宅宅新聞】     蕃Plus+1+1     -->|http://n.yam.com/gamme/otaku/20150618/20150618100277.html|2015-06-18
其他媒体|1878123383|webcars|降价信息|ZHO|2015-06-29 03:33:01|[郑州]  起亚K3S最高现金优惠1.7万元 可试乘试驾|"　　【万车网 郑州行情】近日 万车网郑州站编辑从东风悦达起亚河南新裕隆4S店了解到 购起亚K3S最高现金优惠1.7万元 现车充足 颜色可选 感兴趣的朋友可与经销商联系。具体优惠信息请见下表：　　近期火爆活动：　　【全城最低价 组团买新车】万车网团车活动火爆进行中（点击进入）　起亚K3S郑州地区行情车型指导价（万元）经销商报价（万元）优惠幅度（万元）2014款 1.6L 手动GL10.188.50↘1.682014款 1.6L 自动GL11.189.50↘1.682014款 1.6L 手动GLS11.489.70↘1.682014款 1.6L 自动GLS12.4810.80↘1.682014款 1.6L 自动DLX13.1811.40↘1.682014款 1.6L 自动Premium14.3812.68↘1.702015年6月29日行情 车辆价格随时变动 敬请关注当地市场http://www.webcars.com.cn/万车网制表您询问和购车时说明您是""万车网用户"" 会得到更好的服务！《点击可查看郑州地区起亚4S店》　　与K3不同 起亚K3S前进气格栅尺寸明显缩小 前保险杠采用大嘴式设计 整车设计更加年轻动感。车身尺寸方面 起亚K3S长宽高分别为4365/1780/1460mm 轴距达到2700mm。车身颜色方面 起亚K3S有透明白、钻石银、檀木黑、暗樱红、汉玉白、钛银色和新雅蓝共7款车身颜色可选。【起亚K3S 外观】【起亚K3S 外观】　　内饰方面 起亚K3S与K3整体内饰布局保持高度一致 中控台采用不对称式设计 在搭配黑色仿碳纤维装饰后 车内驾驶氛围凸显运动气息。内饰配色方面 起亚K3S还增加了黑棕配色方案供消费者选择。配置方面 起亚K3S全系标配后扰流板、随速感应自动落锁、带有CD(MP3)+AUX+USB+iPod读取功能的音响系统、前排座椅安全带高度可调、前排电子预紧式安全带等配置。除入门级车型外 余下5款车型均配有倒车雷达。【起亚K3S 内饰】【起亚K3S 内饰】　　动力方面 起亚K3S搭载了1.6L自然吸气发动机 该发动机的最大功率为128马力 峰值扭矩为156N·m。传动方面 与之匹配的是6速手动或6速自动变速箱。　　经销商信息：　　经销商名称：河南新裕隆汽车销售服务有限公司　　经销商地址：郑州市花园北路与开元路交叉口河南汽车贸易中心院内　　经销商电话：0371-65******-*******6　　声明：　　本文中涉及到的车型价格为万车网编辑在经销商处采集到的真实当日价格。由于汽车价格经常变化 并且为单一经销商的个体行为 所以价格仅供参考。具体价格请您致电或到店与经销商详细商谈。文中图片为车型实拍图 价格信息与图片拍摄地点无关。    本文导航         责任编辑：关鑫  关键词：起亚K3S 东风悦达起亚 郑州悦达起亚 起亚k3 福瑞迪 起亚k5 起亚k2 起亚智跑 起亚k3s 起亚狮跑东风悦达起亚 K3S K3 河南新裕隆       查看车型   实时报价  参数配置  实拍图片  热点资讯  评分评论  万车知道"|http://www.webcars.com.cn/review/20150629/109121.html|2015-06-29
其他媒体|1878286407|difang CN|地方频道 > 滚动读报|ZHO|2015-06-29 08:20:02|油价上涨无所惧 k3节能有攻略|今年3月底到5月初期间 国际油价曾发起一波强劲的反弹攻势 国内成品油价格也完成了“三连涨”。汽车用户们开始纷纷寻找一劳永逸的油价破局纾困之道 百公里最低油耗仅6.3升的东风悦达起亚k3由此落入车主眼帘。k3拥有突出的燃油经济性 性价比杰出。其采用起亚先进的1.6升伽马d-cvvt发动机 最大功率可达128马力。同时 1.8升车型采用nud-cvvt发动机 最大功率可达146马力 并无隙配合先进的6速手自一体变速箱 操控随心 淋漓快意。k3最低油耗更可低至百公里仅6.3升 其高性价比在同排量车型里尽享优势。（起亚）|http://difang.gmw.cn/newspaper/2015-06/29/content_107567106.htm|2015-06-29
其他媒体|1878840966|hexun|滚动新闻 > 全部新闻|ZHO|2015-06-29 14:44:02|起亚k3报价及图片 立减3万现金 现车齐全 颜色可选 销售全国|2015款K3秉承“Design KIA”设计理念精髓 在车身前脸和尾部均有全新呈现。前脸全新的前中网颜色 使得虎啸式家族脸谱视觉感受更为动感大气且引人注目。近日 笔者从东风悦达起亚北京金宝龙4S店获悉 目前2015款K3现车充足 颜色可选 全国可售 全系优惠3万元 近期购车综合优惠可达4万 与之前相比优惠大幅增加。欢迎感兴趣的朋友致电详询。　　外地客户可报销两人单程车票！　　近期购车送万元礼包：　　全车膜（进口）、地胶、脚垫、凉垫、把套、麂皮、掸子、发动机护板、车身封釉、地盘封塑、后舱垫、行李架、脚踏板、前后保险杠、DVD导航、原厂导航、倒车影像、倒车雷达、真皮座椅、挡泥板　　销售咨询电话：18001******-*******9508 那经理车型(北京报价)指导价(万)本店店价格(万)价格变化(万)备注1.6L 手动GL2015款10.287.28↓3现车充足1.6L 自动GL2015款11.288.28↓3现车充足1.6L 手动GLS2015款11.488.48↓3现车充足1.6L 自动GLS2015款12.489.48↓3现车充足1.6L 自动DLX2015款13.1810.18↓3现车充足1.6L 自动Premium2015款14.3811.38↓3现车充足1.8L 自动Premium2015款14.9811.98↓3现车充足　　装饰礼包（选装）：　　全车膜（进口）、地胶、脚垫、凉垫、把套、麂皮、掸子、发动机护板、车身封釉、地盘封塑、后舱垫、行李架、脚踏板、前后保险杠、DVD导航、原厂导航、倒车影像、倒车雷达、真皮座椅、挡泥板　　2015款K3车型的前中网颜色变更 后保险杠和排气管也经过了重新设计 DLX AT及以上车型配备了椭圆形的镀铬排气管。2015款K3还新增珍珠白这一可选车身颜色。中控面板位置的空调按钮将增加镀铬装饰 车内还将引入更多软性材料装饰。配置方面 新款K3将全系标配外后视镜加热功能 两款Premium车型都将配备带有加热和通风功能的电动调节前座椅 DLX AT车型则可选装该配置。　　我们秉承“诚信经营 价格合理 双赢合作 服务第一”的服务理念　　更多详情请联系经销商：　　公司名称: 北京金宝龙达汽车4S店　　经营性质: 综合4S店　　联 系 人: 那经理 和我联系　　销售电话: 18001******-*******9508　　公司网址: www.im4s.cn/30875　　公司地址：北京市昌平区北五环立汤路58号　　北京站乘车路线: 北京站-坐2号线地铁到崇文门-转5号线地铁天通苑站下车即到　　北京西站乘车路线: 北京西站-坐9号线地铁到白石桥南-转6号线地铁到东四-转5号线地铁 天通苑站下车即到　　北京南站乘车路线： 北京南站坐4号线地铁到宣武门站-转2号线地铁到崇文门转-5号线地铁 到天通苑站下车即到　　注： 本综合性4S店只为客户提供裸车 仅销往山西 陕西 内蒙古 河南 河北 山东 安徽 甘肃 东北等地 　　联系方式：　　销售电话：18001******-*******8537　　售后电话：***********　　联系人：那经理更多网站功能:汽车大全 汽车报价 汽车资讯网　　如系本站原创文章 转载请注明出处：汽车中国。　　更多汽车新闻关注 请扫码汽车中国公众微信号：（责任编辑：HN666）|http://auto.hexun.com/2015-06-29/177125675.html|2015-06-29
其他媒体|1879238907|hexun|滚动新闻 > 全部新闻|ZHO|2015-06-29 18:31:03|东风起亚k3现车销售优惠高达现金5万元 配置参数安全性能油耗资讯|　　悦达起亚作为起亚在华的合资品牌 K3成为东风悦达起亚旗下引入的第三款K系列车型 K3已经在成都车展亮相 其搭载了与现代朗动相同的动力系统 1.6L及1.8L发动机 并于2012年10月15日左右上市。近日 编辑从北京润通嘉华汽车销售有限公司获悉 东风起亚k3有最新优惠活动 目前该店内东风起亚k3现车销售 面向全国 无限地域 颜色可选 优惠高达现金5万元 购车即赠价值20000万豪华大礼包。对东风起亚k3感兴趣的车友可以联系该店。[联系电话]；*********** 王经理车型(广州报价)指导价(万)4s店价格(万)价格变化(万)备注起亚K3 1.6L MTGL2012款***.***.***.***赠20000万元礼包起亚K3 1.6L ATGL2012款***.***.***.***赠20000元礼包起亚K3 1.6L MTGLS2012款***.***.***.***起亚K3 1.6L ATGLS2012款***.***.***.***起亚K3 1.6L ATDLX2012款13.1810.183.0起亚K3 1.6L ATPremium2012款14.38　　11.383.0　　以上优惠信息为经销商提供 部分价格会与实际情况有差异 真实价格以到店为准 或先致电咨询；*********** 王经理　　东风悦达起亚全新K3相较K2和K5的设计 有了明显区别 十分突出力量感和线条的精炼。在前脸的设计上 采用起亚最高端旗舰车型K9的镀铬直瀑式竖条进气格栅 视觉感受更为大气、稳健；前后大灯都采用LED设计 再配合LED日间行车灯 彰显出浓厚的科技感以及时代感；在精炼线条勾勒下 大倾角前风挡以及溜背式车尾处理都传递出独特的动态肌肉造型美 视觉冲击强烈 让人过目难忘。K3的设计风格 是简约直线美学设计理念的再升华 是对“DESIGN KIA”的完美诠释。　　[推荐商家] 北京润通嘉华汽车销售有限公司[联系电话]*********** 王经理　　[商家地址] 北京市昌平区天通苑北61号　　咨询时若提及是在汽车中国看到的将可享受更多优惠更多网站功能:汽车大全 汽车报价 汽车资讯网　　如系本站原创文章 转载请注明出处：汽车中国。　　更多汽车新闻关注 请扫码汽车中国公众微信号：（责任编辑：HN666）|http://auto.hexun.com/2015-06-29/177132620.html|2015-06-29
其他媒体|1879474847|pconline|论坛-keyword_三星|ZHO|2015-06-29 21:08:01|一大堆小东西 喜欢的来秒！|欧特斯 卡通创意可爱叮当猫16G迷你优盘包邮高速优盘个性定制礼品【今日特价秒杀19.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/HPNEG1y 游戏有线USB办公键盘CFLOL 电脑笔记本台式键盘 防水超薄静音包邮【今日特价秒杀17.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/dkHEG1y 鼎铃正品电动男用鼻毛修剪器刮鼻毛器剃鼻毛充电鼻毛修剪特价包邮【今日特价秒杀15.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/qCFEG1y B-LINK 四天线无线路由器穿墙王 家用宽带智能无限WIFI发射ap迷你【今日特价秒杀59.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/7lIEG1y 宏邦蒸脸迷你挂烫机手持熨烫机电熨斗蒸汽美容家用小型便携式旅行【今日特价秒杀29.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/ClJEG1y B-LINK USB无线网卡 迷你WIFI接收发射器手机台式机电脑笔记本AP【今日特价秒杀19.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/JBHEG1y 超界电子称体重秤家用电子秤称精准人体秤健康秤体重计智能称包邮【今日特价秒杀39.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/99GEG1y ione/艾旺 PA-101 酸奶机全自动 家用不锈钢胆多功能恒温正品特价【今日特价秒杀19.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/AbDEG1y 十全十美 Q20B蓝牙多媒体2.1低音炮音响有源笔记本台式电脑小音箱【今日特价秒杀128.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/16DEG1y X·AI A3无线蓝牙手机免提迷你插卡小音箱金属创意便携低音炮音响【今日特价秒杀29.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/UZDEG1y 多功能鸡蛋杯卷蛋器卷蛋机早餐机蒸蛋器煮蛋器家用懒人早餐神器【今日特价秒杀29.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/k3EEG1y 思考个性迷你小精灵u盘16g创意女生礼品高速车载优盘16g特价免邮【今日特价秒杀19.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/vx8EG1y ZTE/中兴 小球音箱便携式迷你小音响小米魅族苹果手机扩音器通用【今日特价秒杀35.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/o2GEG1y 梦族平板支架床头床上夹子懒人苹果mini架子电脑手机通用ipad支架【今日特价秒杀18.80元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/Rq5EG1y SAST/先科 mx-505蓝牙音箱 电脑手机迷你插卡小音响低音炮收音机【今日特价秒杀45.01元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/Qf9EG1y 拓普赛特 K16四核网络机顶盒wifi无线高清硬盘播放器电视机顶盒子【今日特价秒杀299.03元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/TG4EG1y FS372飞科剃须刀男士电动刮胡刀充电式剃胡须刀全身水洗须刨正品【今日特价秒杀99.02元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/RZ8EG1y 朗威Rs831电动剃须刀电动双头充电式刮胡刀男剃胡刀胡须正品特价【今日特价秒杀25.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/KH9EG1y 飞科剃须刀FS360男士飞科电动剃须刀刮胡刀充电式胡须刀正品包邮【今日特价秒杀65.01元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/OO4EG1y 上海红心电熨斗RH183家用 蒸汽熨斗 手持挂式迷你电烫斗正品包邮【今日特价秒杀57.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/5C7EG1y 买二有礼 手提电脑包A4文件包多功能收纳包 办公学习用品【今日特价秒杀9.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/0guDG1y 第一眼 HP990木质USB2.0低音炮手机笔记本台式迷你电脑音响小音箱【今日特价秒杀19.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/ZGzDG1y 真汉子RSCF-8237双头电动剃须刀刮胡刀充电式浮动胡须刀水洗刀头【今日特价秒杀19.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/mG2EG1y 中兴 原装重低音小米魅族三星通用带麦线控有线耳机耳塞式入耳式【今日特价秒杀79.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/tF1EG1y 中兴无线手机蓝牙音响电脑平板迷你音箱便携式低音炮立体声户外【今日特价秒杀69.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/lrvDG1y ZTE/中兴 T630 商务蓝牙耳塞挂耳式耳机4.0小米三星苹果4.1通用【今日特价秒杀68.80元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/61sDG1y 中兴青花瓷移动电源通用毫安手机超薄迷你聚合物充电宝充电宝【今日特价秒杀68.80元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/uJuDG1y ZTE中兴手机通用充电器USB直充直冲插头套装旅行车载套装zte安卓【今日特价秒杀59.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/OksDG1y 飞科电吹风大功率家用吹风机学生旅游冷热风电吹风机宿舍FH6622【今日特价秒杀49.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/xVvDG1y 飞科成人通用理发器充电式剃头刀电推剪儿童剃发套装电剪推头剪发【今日特价秒杀69.01元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/xCiDG1y 女士专用脱毛器充电动剃毛器男女用刮毛刀腋下私处剃腋毛阴毛腿毛【今日特价秒杀55.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/8RkDG1y 飞科理发器电动推剪头发成人儿童电推子充电式剃发剃头刀家用专业【今日特价秒杀59.01元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/gOmDG1y   评分  分享|http://itbbs.pconline.com.cn/es/52343490.html|2015-06-29
其他媒体|1879474848|pconline|论坛-keyword_三星|ZHO|2015-06-29 21:08:01|【特价数码家电】正品行货 秒到赚到！|欧特斯 卡通创意可爱叮当猫16G迷你优盘包邮高速优盘个性定制礼品【今日特价秒杀19.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/HPNEG1y 游戏有线USB办公键盘CFLOL 电脑笔记本台式键盘 防水超薄静音包邮【今日特价秒杀17.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/dkHEG1y 鼎铃正品电动男用鼻毛修剪器刮鼻毛器剃鼻毛充电鼻毛修剪特价包邮【今日特价秒杀15.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/qCFEG1y B-LINK 四天线无线路由器穿墙王 家用宽带智能无限WIFI发射ap迷你【今日特价秒杀59.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/7lIEG1y 宏邦蒸脸迷你挂烫机手持熨烫机电熨斗蒸汽美容家用小型便携式旅行【今日特价秒杀29.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/ClJEG1y B-LINK USB无线网卡 迷你WIFI接收发射器手机台式机电脑笔记本AP【今日特价秒杀19.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/JBHEG1y 超界电子称体重秤家用电子秤称精准人体秤健康秤体重计智能称包邮【今日特价秒杀39.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/99GEG1y ione/艾旺 PA-101 酸奶机全自动 家用不锈钢胆多功能恒温正品特价【今日特价秒杀19.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/AbDEG1y 十全十美 Q20B蓝牙多媒体2.1低音炮音响有源笔记本台式电脑小音箱【今日特价秒杀128.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/16DEG1y X·AI A3无线蓝牙手机免提迷你插卡小音箱金属创意便携低音炮音响【今日特价秒杀29.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/UZDEG1y 多功能鸡蛋杯卷蛋器卷蛋机早餐机蒸蛋器煮蛋器家用懒人早餐神器【今日特价秒杀29.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/k3EEG1y 思考个性迷你小精灵u盘16g创意女生礼品高速车载优盘16g特价免邮【今日特价秒杀19.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/vx8EG1y ZTE/中兴 小球音箱便携式迷你小音响小米魅族苹果手机扩音器通用【今日特价秒杀35.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/o2GEG1y 梦族平板支架床头床上夹子懒人苹果mini架子电脑手机通用ipad支架【今日特价秒杀18.80元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/Rq5EG1y SAST/先科 mx-505蓝牙音箱 电脑手机迷你插卡小音响低音炮收音机【今日特价秒杀45.01元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/Qf9EG1y 拓普赛特 K16四核网络机顶盒wifi无线高清硬盘播放器电视机顶盒子【今日特价秒杀299.03元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/TG4EG1y FS372飞科剃须刀男士电动刮胡刀充电式剃胡须刀全身水洗须刨正品【今日特价秒杀99.02元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/RZ8EG1y 朗威Rs831电动剃须刀电动双头充电式刮胡刀男剃胡刀胡须正品特价【今日特价秒杀25.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/KH9EG1y 飞科剃须刀FS360男士飞科电动剃须刀刮胡刀充电式胡须刀正品包邮【今日特价秒杀65.01元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/OO4EG1y 上海红心电熨斗RH183家用 蒸汽熨斗 手持挂式迷你电烫斗正品包邮【今日特价秒杀57.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/5C7EG1y 买二有礼 手提电脑包A4文件包多功能收纳包 办公学习用品【今日特价秒杀9.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/0guDG1y 第一眼 HP990木质USB2.0低音炮手机笔记本台式迷你电脑音响小音箱【今日特价秒杀19.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/ZGzDG1y 真汉子RSCF-8237双头电动剃须刀刮胡刀充电式浮动胡须刀水洗刀头【今日特价秒杀19.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/mG2EG1y 中兴 原装重低音小米魅族三星通用带麦线控有线耳机耳塞式入耳式【今日特价秒杀79.90元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/tF1EG1y 中兴无线手机蓝牙音响电脑平板迷你音箱便携式低音炮立体声户外【今日特价秒杀69.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/lrvDG1y ZTE/中兴 T630 商务蓝牙耳塞挂耳式耳机4.0小米三星苹果4.1通用【今日特价秒杀68.80元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/61sDG1y 中兴青花瓷移动电源通用毫安手机超薄迷你聚合物充电宝充电宝【今日特价秒杀68.80元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/uJuDG1y ZTE中兴手机通用充电器USB直充直冲插头套装旅行车载套装zte安卓【今日特价秒杀59.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/OksDG1y 飞科电吹风大功率家用吹风机学生旅游冷热风电吹风机宿舍FH6622【今日特价秒杀49.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/xVvDG1y 飞科成人通用理发器充电式剃头刀电推剪儿童剃发套装电剪推头剪发【今日特价秒杀69.01元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/xCiDG1y 女士专用脱毛器充电动剃毛器男女用刮毛刀腋下私处剃腋毛阴毛腿毛【今日特价秒杀55.00元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/8RkDG1y 飞科理发器电动推剪头发成人儿童电推子充电式剃发剃头刀家用专业【今日特价秒杀59.01元包邮】【淘宝链接 复制打开】http://s.click.taobao.com/gOmDG1y   评分  分享|http://itbbs.pconline.com.cn/es/52343492.html|2015-06-29
其他媒体|1886285305|hefei|合肥专区|ZHO|2015-07-03 12:51:01|2015年日语二级考试 答案《★*********★》|"2015年日语二级考试 答案《★*********★》  2015年日语二级考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年日语二级考试真题答案-2015年日语二级试题及 答案-2015年日语二级考试时间-2015年日语二级考试科目-2015年日语二级考试大纲-2015年日语二级考前答案-2015年日语二级答案【Q*********包过】-2015年日语二级考试资料【Q*********包过】-2015年日语二级复习资料-2015年日语二级考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级日语二级著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年日语二级考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级日语二级考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年日语二级考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级日语二级 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年日语二级考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年日语二级考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级日语二级考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级日语二级考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级日语二级考试 答案=*********.祈福2015年日语二级考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年日语二级考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年日语二级考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级日语二级考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年日语二级考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级日语二级考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年日语二级考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年日语二级考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年日语二级考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年日语二级考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年日语二级考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年日语二级考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级日语二级考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级日语二级答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级日语二级考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年日语二级考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年日语二级考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年日语二级考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年日语二级考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级日语二级考试英语考式考式 考式 答案= 高级高级日语二级考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年日语二级考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年日语二级考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年日语二级考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年日语二级考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级日语二级答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级日语二级 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年日语二级考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级日语二级考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年日语二级考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级日语二级考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年日语二级考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级日语二级考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年日语二级考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级日语二级考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年日语二级考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年日语二级考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年日语二级考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15307954&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-07-03
其他媒体|1886305882|hefei|合肥专区|ZHO|2015-07-03 13:06:01|2015年日语等级N1考试 答案《★********★》|"2015年日语等级N1考试 答案《★********★》  2015年日语等级N1考试 答案【通过率100%卡卡客服Ｑ********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年日语等级N1考试真题答案-2015年日语等级N1试题及 答案-2015年日语等级N1考试时间-2015年日语等级N1考试科目-2015年日语等级N1考试大纲-2015年云南丽江市属事业单位招聘考前答案-2015年日语等级N1答案【Q********包过】-2015年日语等级N1考试资料【Q********包过】-2015年日语等级N1复习资料-2015年云南丽江市属事业单位招聘考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级河南省考著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年日语等级N1考试 答案=********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级河南省考考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @' }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年日语等级N1考试 答案 试题 真题 时间 科目〃Ｑ******** ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年日语等级N1考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年日语等级N1考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级河南省考考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级河南省考考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级河南省考考试 答案=********.祈福2015年云南丽江市属事业单位招聘考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年日语等级N1考试 考式 答案=********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年日语等级N1考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=********人时简累 会受苦 正高级高级河南省考考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =********.祈福2015年日语等级N1考试 考式 答案=********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级河南省考考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=********.祈福2015年日语等级N1考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=******** ^1 q) ~# t: {/ h/ J【=********.祈福2015年日语等级N1考试 考式 答案=******** W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年日语等级N1考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. ********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年日语等级N1考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=********.祈福2015年日语等级N1考试 考式 答案=********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级河南省考考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级河南省考答案【Q********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级河南省考考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=******** 2015年日语等级N1考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年日语等级N1考试 考式 答案=********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年日语等级N1考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=******** 2015年日语等级N1考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级河南省考考试英语考式考式 考式 答案= 高级高级河南省考考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W********=******** 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^ ********_100%】哪个2015年日语等级N1考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年日语等级N1考试 考式 答案=********.+ F; ~ C( X7 G$ ?$ I祈福2015年日语等级N1考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年日语等级N1考试 考式 答案=********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级河南省考答案【Q********】9 I' [+ v* p3 m' Q =********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级河南省考 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年日语等级N1考试 考式 答案=********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级河南省考考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年日语等级N1考试 考式 答案=********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级河南省考考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”********.祈福2015年日语等级N1考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级河南省考考试/ J7 J' y9 ]5 c5 w; D答案=********.祈福2015年日语等级N1考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级河南省考考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年日语等级N1考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案********.祈福2015年云南丽江市属事业单位招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年日语等级N1考试 答案Ｑ********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15308003&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-07-03
其他媒体|1886324660|hefei|合肥专区|ZHO|2015-07-03 13:19:02|2015年日语三级考试 答案《★*********★》|"2015年日语三级考试 答案《★*********★》  2015年日语三级考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年日语三级考试真题答案-2015年日语三级试题及 答案-2015年日语三级考试时间-2015年日语三级考试科目-2015年日语三级考试大纲-2015年日语三级考前答案-2015年日语三级答案【Q*********包过】-2015年日语三级考试资料【Q*********包过】-2015年日语三级复习资料-2015年日语三级考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级日语三级著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年日语三级考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级日语三级考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年日语三级考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级日语三级 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年日语三级考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年日语三级考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级日语三级考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级日语三级考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级日语三级考试 答案=*********.祈福2015年日语三级考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年日语三级考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年日语三级考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级日语三级考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年日语三级考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级日语三级考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年日语三级考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年日语三级考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年日语三级考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年日语三级考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年日语三级考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年日语三级考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级日语三级考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级日语三级答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级日语三级考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年日语三级考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年日语三级考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年日语三级考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年日语三级考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级日语三级考试英语考式考式 考式 答案= 高级高级日语三级考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年日语三级考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年日语三级考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年日语三级考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年日语三级考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级日语三级答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级日语三级 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年日语三级考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级日语三级考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年日语三级考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级日语三级考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年日语三级考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级日语三级考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年日语三级考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级日语三级考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年日语三级考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年日语三级考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年日语三级考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15308087&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-07-03
기타|1886745420|ngzb|新闻互动|ZHO|2015-07-03 17:45:01|银联国际在韩持续发力 创新服务提升用卡体验|"马上注册 结交更多好友 享用更多功能 让你轻松玩转南宁您需要 登录 才可以下载或查看 没有帐号？立即注册  x银联国际在韩持续发力 创新服务提升用卡体验8 h( a0 n' e7 G& q3 M　　记者7月3日最新获悉 银联国际已在韩国推出退税即时到账服务 并与主流机构合作发行当地首张银联“闪付”卡 还在商户受理环境优化、丰富用卡权益等多个领域取得新进展。+ c2 C- A0 P1 N4 w' Z: n| k$ W- b8 k  T2 Z/ T. b& _( n+ Z) ?' {* t"" F　　在韩国旅游业受MERS疫情影响的背景下 银联国际致力于在淡季不断提升创新能力和服务水平 支持韩国政府振兴当地经济和旅游业发展。近期 银联国际在明洞、江南、梨泰院等首尔主要观光区检查 以进一步优化受理质量 确保MERS疫情缓解后 游客再次大量涌入韩国时可以享受更优质的银联卡支付服务。5 A+ [8 P' H| M"" j1 P: M| R3 g3 @| M7 F; E( v7 n　　推出退税即时到账服务+ U  f6 ?| l7 s"" J' w| V+ x( Z0 m- ^; A　　银联国际与韩国最大的退税服务公司Global Tax Free（GTF）合作 首次推出中国境内银联卡（卡号以62开头）持卡人在韩退税即时到账服务 这也是迄今为止当地最快捷的退税服务 标志着韩国的银联卡产品和服务创新又获新进展。3 P0 m4 r. Q9 Q7 x2 `4 t; s( M1 a1 F% S# V　　游客在GTF特约商户购物后 可在市内退税服务台领取退税单 离境时在各大机场和港口海关盖章后 向GTF退税窗口提供姓名、护照号、国籍、银联卡卡号和身份证后6位 即可申请退税 税款即时返还至该银联卡中。  w# h( k/ `% C4 i: T6 C- U% E5 @3 z0 }6 d3 P　　创新支付提升用卡体验1 X| T"" {9 _4 c5 g2 K6 t: m3 T) T3 ^3 w- u& ?　　再次扩大银联“闪付”服务范围。近期 韩国受理银联“闪付”卡的范围进一步扩大。银联卡持卡人已可在首尔东大门斗塔购物中心及8100余家GS25便利店体验快捷、便利、安全的“拍”卡支付。更多便利店、免税店、咖啡厅等将陆续开通。: `( q3 k+ n* k3 }4 @$ O* @/ e/ i- X3 P  M* o　　本周 银联国际还与韩国主流机构正式合作 发行首张针对韩国人的银联“闪付”卡 近期还将在移动端推出非接产品 支持本地居民在全球500多万台“闪付”终端“拍”卡支付。0 s& L) \) v) \+ q* Y$ u: i2 z9 X/ u5 o$ B; W+ V1 C+ [　　携手T-money创新交通支付。为了解决游客赴韩后购买韩国T-Money交通卡的不便 银联国际还与韩国智能卡公司合作 9月中旬开始 中国境内银联“闪付”卡持卡人便可通过手机 在韩国使用T-Money交通卡的服务。此举为即将到来的国庆出游高峰提供了更便利的解决方案。/ r7 W(  0 E4 q% O' N5 v$ }* e( w2 X1 N9 l4 [　　启动6万韩国网上商户大型优惠: U| U) j% ~"" m1 [) ]- n- Z; R9 }3 f+ R: p　　在访韩游客大幅减少的情况下 银联国际7月将启动韩国网上商户大型优惠活动 让银联卡持卡人不出国门也能买到心仪的韩国商品。目前 韩国已有6万多家网上商户可用银联卡支付 包括Lotte.com、Gmarket、新罗免税店等知名线上商户 这一范围还在不断扩大。+ @6 T) C6 n6 y  d) P| n1 l( ~| z　　提升韩国持卡人出行支付体验8 a. u4  2 Y1 ~) S/ L% y$ V"" X) C' j' b( g) b& g4 @　　随着当地银联卡产品和权益体系的不断丰富 韩国居民对银联品牌也日益认可 现在每5个韩国人就拥有一张银联卡。今年 银联国际携手友利卡公司发行了“友利自由旅行卡” 该卡在韩国人最喜欢的亚洲五国提供多项旅游相关优惠礼遇 包括机票九折、免费使用银联休息室、热门景点八五折优惠、乐天免税店VIP金卡升级等 吸引了众多韩国人办卡。"" q1 j; t8 }0 Y1 q0 m( H. T( c* u& s  C' c. Z( E"" t　　与全球其他银联卡持卡人一样 韩国持卡人也可在仁川机场享受直通列车特价票、机场免税店最高6万元折扣、仁川银联咖啡厅免费上网及免费咖啡礼遇 并在日本、香港、美国等地多个热门旅游目的地享受丰富优惠及权益。' [* a9 T. {' ]""  ( \"" _0 X' a4 V"" {) U& u* ]  ^+ W　　目前 几乎所有韩国签名受理商户都接受银联信用卡 近120万家商户可用银联卡进行密码支付 几乎所有出租车都可以刷银联信用卡支付。$ l; F0 a6 U9 s| T"" H: e! z: U- G9  % z7 Z- c| t　　关于银联国际: `9 u$ [8 B$ B% O) m3 b; e. }5 z1 g% s+ ^* s　　银联国际是中国银联负责运营国际业务的子公司 以会员制吸引全球合作伙伴 拓展银联卡境外受理网络 扩大银联卡发行和使用 开展创新支付的跨境应用 提升银联品牌的国际影响力。通过与全球300多家机构合作 目前银联境外受理网络已延伸到150个国家和地区 40个国家和地区发行了银联卡。银联国际正在为全球最大的持卡人群提供优质、高效、安全的跨境支付服务 并为越来越多境外银联卡持卡人提供日益便利的本地化服务。/ R5 p"" W  _( k% h9 B1 Q7 A6 n1 G2 T8 L/ z% N$ @- {6 s　　如欲了解银联国际更多信息 请访问：www.unionpayintl.com 或关注“银联国际”新浪微博、“银联国际”微信公众号 下载“银联国际”手机APP。; ^! T1 S8 t! E$ W| K7 ^  G) n# o6 H! s& \0 C' ^- M　　媒体联系：*****@************.***' }% d1 r1 U| \7 r/ @! _* @% g& D"" }"" a"" U; M"" q/ c　　登录/注册后可看大图图片2.jpg (30.26 KB| 下载次数: 0)下载附件 保存到相册10 分钟前 上传</ignore_js_op>- X+ b+ K  c/ m2 r4 e! r9 ~! z2 ?8 U# p7 f/ z3 z$ C*  & I) {9 t　　　APP中文版                  APP英文版                   微信服务号                  微信订阅号/ d6 T$ J/ q  M2 S& r% L"" \2 Q) k5 V| s$ M4 `3 k3 F9 f2 s; ?| D韩国政府| 身份证| 服务公司| 旅游业| 服务台"|http://www.ngzb.com.cn/forum.php?mod=viewthread&tid=946280&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline|2015-07-03
其他媒体|1892378563|hefei|合肥专区|ZHO|2015-07-07 10:25:02|2015年甘肃一万名考试 答案《★*********★》|"2015年甘肃一万名考试 答案《★*********★》  2015年甘肃一万名考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年甘肃一万名考试真题答案-2015年甘肃一万名试题及 答案-2015年甘肃一万名考试时间-2015年甘肃一万名进村进社考试科目-2015年甘肃一万名考试大纲-2015年甘肃一万名考前答案-2015年甘肃一万名答案【Q*********包过】-2015年甘肃一万名考试资料【Q*********包过】-2015年甘肃一万名复习资料-2015年甘肃一万名考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级甘肃一万名著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年甘肃一万名考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级甘肃一万名考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年甘肃一万名考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年甘肃一万名考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年甘肃一万名考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级甘肃一万名考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级甘肃一万名考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级甘肃一万名考试 答案=*********.祈福2015年甘肃一万名进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年甘肃一万名考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年甘肃一万名考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级甘肃一万名考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年甘肃一万名考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级甘肃一万名考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年甘肃一万名考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年甘肃一万名考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年甘肃一万名考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年甘肃一万名考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年甘肃一万名考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级甘肃一万名考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级甘肃一万名答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级甘肃一万名考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年甘肃一万名考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年甘肃一万名考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年甘肃一万名考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年甘肃一万名考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级甘肃一万名考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年甘肃一万名考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年甘肃一万名考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年甘肃一万名考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年甘肃一万名考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级甘肃一万名答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级甘肃一万名 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年甘肃一万名考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级甘肃一万名考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年甘肃一万名考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级甘肃一万名考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年甘肃一万名考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级甘肃一万名考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年甘肃一万名考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级甘肃一万名考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年甘肃一万名考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年甘肃一万名考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15316846&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-07-07
其他媒体|1892425014|hefei|合肥专区|ZHO|2015-07-07 10:55:01|2015年甘肃10000名考试 答案《★*********★》|"2015年甘肃10000名考试 答案《★*********★》  2015年甘肃10000名考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年甘肃10000名考试真题答案-2015年甘肃10000名试题及 答案-2015年甘肃10000名考试时间-2015年甘肃10000名进村进社考试科目-2015年甘肃10000名考试大纲-2015年甘肃10000名考前答案-2015年甘肃10000名答案【Q*********包过】-2015年甘肃10000名考试资料【Q*********包过】-2015年甘肃10000名复习资料-2015年甘肃10000名考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级甘肃10000名著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年甘肃10000名考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级甘肃10000名考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年甘肃10000名考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年甘肃10000名考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年甘肃10000名考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级甘肃10000名考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级甘肃10000名考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级甘肃10000名考试 答案=*********.祈福2015年甘肃10000名进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年甘肃10000名考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年甘肃10000名考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级甘肃10000名考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年甘肃10000名考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级甘肃10000名考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年甘肃10000名考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年甘肃10000名考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年甘肃10000名考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年甘肃10000名考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年甘肃10000名考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级甘肃10000名考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级甘肃10000名答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级甘肃10000名考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年甘肃10000名考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年甘肃10000名考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年甘肃10000名考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年甘肃10000名考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级甘肃10000名考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年甘肃10000名考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年甘肃10000名考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年甘肃10000名考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年甘肃10000名考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级甘肃10000名答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级甘肃10000名 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年甘肃10000名考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级甘肃10000名考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年甘肃10000名考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级甘肃10000名考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年甘肃10000名考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级甘肃10000名考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年甘肃10000名考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级甘肃10000名考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年甘肃10000名考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年甘肃10000名考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15316898&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-07-07
其他媒体|1893343269|zhidao_baidu|生活|ZHO|2015-07-07 20:04:02|东风悦达起亚k3gls有几个颜色|来自：手机知道江苏|http://zhidao.baidu.com/question/1767937012529940540.html?entry=qb_browse_default|2015-07-07
其他媒体|1893977081|webcars|降价信息|ZHO|2015-07-08 04:01:03|[郑州]  东风悦达起亚K3S最高现金优惠1.7万元|"　　【万车网 郑州行情】近日 万车网郑州站编辑从东风悦达起亚河南新裕隆4S店了解到 购起亚K3S最高现金优惠1.7万元 现车充足 颜色可选 感兴趣的朋友可与经销商联系。具体优惠信息请见下表：　　近期火爆活动：　　【全城最低价 组团买新车】万车网团车活动火爆进行中（点击进入）　起亚K3S郑州地区行情车型指导价（万元）经销商报价（万元）优惠幅度（万元）2014款 1.6L 手动GL10.188.60↘1.582014款 1.6L 自动GL11.189.50↘1.682014款 1.6L 手动GLS11.489.78↘1.702014款 1.6L 自动GLS12.4810.78↘1.702014款 1.6L 自动DLX13.1811.48↘1.702014款 1.6L 自动Premium14.3812.68↘1.702015年7月8日行情 车辆价格随时变动 敬请关注当地市场http://www.webcars.com.cn/万车网制表您询问和购车时说明您是""万车网用户"" 会得到更好的服务！《点击可查看郑州地区起亚4S店》　　与K3不同 起亚K3S前进气格栅尺寸明显缩小 前保险杠采用大嘴式设计 整车设计更加年轻动感。车身尺寸方面 起亚K3S长宽高分别为4365/1780/1460mm 轴距达到2700mm。车身颜色方面 起亚K3S有透明白、钻石银、檀木黑、暗樱红、汉玉白、钛银色和新雅蓝共7款车身颜色可选。【起亚K3S 外观】【起亚K3S 外观】　　内饰方面 起亚K3S与K3整体内饰布局保持高度一致 中控台采用不对称式设计 在搭配黑色仿碳纤维装饰后 车内驾驶氛围凸显运动气息。内饰配色方面 起亚K3S还增加了黑棕配色方案供消费者选择。配置方面 起亚K3S全系标配后扰流板、随速感应自动落锁、带有CD(MP3)+AUX+USB+iPod读取功能的音响系统、前排座椅安全带高度可调、前排电子预紧式安全带等配置。除入门级车型外 余下5款车型均配有倒车雷达。【起亚K3S 内饰】【起亚K3S 内饰】　　动力方面 起亚K3S搭载了1.6L自然吸气发动机 该发动机的最大功率为128马力 峰值扭矩为156N·m。传动方面 与之匹配的是6速手动或6速自动变速箱。　　经销商信息：　　经销商名称：河南新裕隆汽车销售服务有限公司　　经销商地址：郑州市花园北路与开元路交叉口河南汽车贸易中心院内　　经销商电话：0371-65******-*******6　　声明：　　本文中涉及到的车型价格为万车网编辑在经销商处采集到的真实当日价格。由于汽车价格经常变化 并且为单一经销商的个体行为 所以价格仅供参考。具体价格请您致电或到店与经销商详细商谈。文中图片为车型实拍图 价格信息与图片拍摄地点无关。    本文导航         责任编辑：关鑫  关键词：起亚K3S 东风悦达起亚 郑州悦达起亚 起亚k3 福瑞迪 起亚k5 起亚k2 起亚智跑 起亚k3s 起亚狮跑东风悦达起亚 K3S K3 河南新裕隆       查看车型   实时报价  参数配置  实拍图片  热点资讯  评分评论  万车知道"|http://www.webcars.com.cn/review/20150708/109351.html|2015-07-08
기타|1894408882|xda|三星Galaxy S III I9308 RSS|ZHO|2015-07-08 11:22:02|2015年甘肃10000名考试 真题%答-案【+15609+6705】过关*付 2015年甘肃10000名考前时间及试题资...|"[游戏分享]2015年甘肃10000名考试 真题%答-案【+15609+6705】过关*付 2015年甘肃10000名考前时间及试题资...[复制链接]  **************当前在线UID*******阅读权限10好友0帖子4精华0积分1注册时间2015-7-8最后登录2015-7-8门户文章0 精华0帖子4积分1 汉堡9 个注册时间2015-7-8发消息 发表于 1 分钟前 显示全部楼层 阅读模式 注册个账号还能参加论坛各种活动哦~您需要 登录 才可以下载或查看 没有帐号？立即注册  x2015年甘肃10000名考试 真题%答-案【+15609+6705】过关*付+ v' T| m1 N1 u3 L& k: y2015年甘肃10000名考前时间及试题资料+卡卡********** V4; \0 T6 ?: _9 X4 Z  i2 c7 G5 \% q* R4 D4 c! B; j8 v1 a* _. e2015年甘肃10000名考试【真题】+2015年甘肃10000名考前时间及试题资料+***.***.***.***.***.***.***.***.5.(通过率100%)壹手打造.100%保证选 择我们=选 择成 功原题操作[诚信第一| 效率第一|考试大纲、考试真题、考试科目、考试资料4 ~"" E% a1 c& ~% w2 d- l6 q| A3 D2 o( @  G5 t# R1 g7 O0 W  `) Y6 {: z"" I/ W* u' f【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】'  / p( \"" x7 y6 f/ w+ e$ Y. l$ n# t【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】* c. y' x& ]4 d* m. A& p/ ]6 l: D4 o6 p* {% M' d9 p9 q& t/ z; s| C5 D& q  f3 q0 L: I2 M( ]9 [2 }# s# U6 x- ]"" J+ F# M5 e服   ~' r1 i% w3 L$ m4 n4 m"" d% ?"" Y/ Z4 R& y【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】| @5 D; w9 G4 e% Y; r# Z"" z* U2 g$ d; A5 G4 i* N* P( I- ~! V- Y- z0 q6 q9 e1 m| R服 # H4 [5 R% z# D6 Q: S1 W# w9 K| l  o& U& E2 O; q- ?4 V! _/ b& [( Y% O- m6 D【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】 【+***.***.***.***.***.***.***.***.5.】6 m"" l"" B' A4 Z0 E. }6 Q( r) B$ Q6 N$ {1 Z# j/ G: z* I( l% L2 N) k3 s服 ' M. g(  9 g# Y9 U5 s"" D! p# M+ e8 T- a' ~' W; H# d9 s& t8 F8 Q$ f2015年甘肃10000名考试卷答题+「***.***.***.***.***.***.***.***.5.」& M6 ~9 Y6 n$ Y8 V# t) Q3 d0 \. Y  A# ]* [0 {9 t- v( ?7 s* h0 p; y4 U+ n7 N* [+ M( L  j6 R 2015年甘肃10000名考前时间及试题资料+***.***.***.***.***.***.***.***.5.(通过率100%)壹手打造.100%保证选 择我们=选 择成 功原题操作[诚信第一| 效率第一|考试大纲、考试真题、考试科目、考试资料8 M& R. e% ^2 C. s) P- ?2 Y: \$ S9 j) @% F) R8 O 2015年甘肃10000名考前时间及试题资料+***.***.***.***.***.***.***.***.5.考前试题有个小和尚 每天早上负责清扫寺庙院子里的落叶。清晨起床扫落叶实在是一件苦差事 尤其在秋冬之际 每一次起风时 树叶总随风飞舞落下。+***.***.***.***.***.***.***.***.5. +***.***.***.***.***.***.***.***.5. +***.***.***.***.***.***.***.***.5. +***.***.***.***.***.***.***.***.5.& T$ ~. l* j- f! {9 o"" R每天早上都需要花费许多时间才能清扫完树叶 这让小和尚头痛不已。他一直想要找个好办法让自己轻松些。后来有个和尚跟他说：“你在明天打扫之前先用力摇树 把落叶统统摇下来 后天就可以不用扫落叶了。”$ Z. ^# M8 y* B6 t6 w* Q0 E; E% C"" i9 R* L# s5 y) N3 Q/ ~* Y; \+ e% i) J3 k6 f1 r. p! Q7 m; t7 K8 U& X0 O& p) }* \' g: L* n$ `. r1 c4 i; K; K+ e8 n3 d; J! k3 x1 \# v1 A& p 6 z"" z- l- M* u# ]$ {     ^* c& c' K| e3 v/ ^# v' I9 v+ g7 j1 @7 }0 j$ I. S1 j0 L; w! t& l) h小和尚觉得这是个好办法 于是隔天他起了个大早 使劲地猛摇树干 这样他就可以把今天跟明天的落叶一次扫干净了。一整天小和尚都非常开心。+ Q3 Z2 U6 N; F+ @* S8 A! U7 R+ B1 f. O4 X$ M% a9 C| z/ `. c9 i| n* P' o+ s3 o8 U7 d; ^: R- g3 r. x1 J  l3 C5 `| U- a2 o0 G$ H4 K2 v  H; P$ U3 i! e6 A% Z; [+ ^5 b% N% A# i( H"" H6 @- Y! T) p+ x* g 1 S. k7 v1 U: A' {第二天 小和尚到院子一看 不禁傻眼了 院子里如往日一样落叶满地。9 K/ I"" d: `2 Z9 `- C: H7 _* ]+ R) }. x0 d/ G8 \! ]$ q1 u. m* n; f# N9 ?4 z: @$ F7 }5 b4 V8 i$ k; A2 n! ^2 d+ N7 A5 l* _/ V. Y. V& w& z: F0 r7 l7 U"" W4 u3 Y: n# q8 U& n这时老和尚走了过来 对小和尚说：“傻孩子 无论你今天怎么用力 明天的落叶还是会飘下来。”小和尚终于明白了 世上有很多事是无法提前的 惟有认真地活好当下 才是最真实的人生态度。青山遮不住 毕竟东流去。该发生的你怎么阻挡也阻挡不了 不会发生的你再努力也没有用。把当下的事情做好了 就无怨无悔。9 ~% D$ X6 I( P| J; A5 W! D3 O& X* y+ A"" g"" d: x"" X4 ]( F0 [( `* z' d% l( \# K9 q! L9 z; [$ k1 t# }: A& m; d5 l0 [6 @6 n. f' ]; E1 M: n' }8 Z7 S2 S/ {' B: M- d$ X( P生活原本没有痛苦- S9 j. e8 W& g: J| E% h. I! ^7 h+ G8 K' ?| O9 m- u1 Y+ ^! L8 u* o$ P$ F"" `: H+ x1 w! B' j7 Y6 f& N( ]. J. r% U4 e* Q. X! s  s  K. k) V5 B* t9 I 0 v2 b- S# n; A8 ?6 Y. e  ^* f6  ! E+ H7 ]/ l& I3 n: Q) ~  l3 {0 _| }- I8 Z生活原本没有烦恼 当欲望之火被点燃后 烦恼就来敲你的心门了。* V* h( W/ f$ i* i. `; w. D6 s5 f. s0 R- h7 m"" P5 R' L. G- C"" D* M6 X( s"" u; o) k8 ^9 B"" q!  : o( F7 N# f7 R1 q% M& Z4 e1 @( y2 I(  . Z0 V( G1 K2 K ) u* r+ K7 Q| u3 P  d/ C. z# h- T6 n; i0 B* H& g* A! X: I8 g7 R| C生活原本没有痛苦 当你开始计较得失 贪求更多时 痛苦便来缠身了。+ k| a% f9 ]2 E8 }( n2 M9 u$ E! A+ e"" O& R0 A9 m| K. c$ B- r. F8 e2 K"" m' i# n$ A3 z5 Z' d9 m& ^1 l9 g: W( c& j& W+ a& Q+ C1 O# }- d' k7 T: @# i! J* U' N/ V. M  ^; r) _) `  \8 e( M : g1 b* q& O# _/ K6 D$ t/ a"" }- H2 i: {: P5 N: a% f0 E7 v; o1 ~3 ?; z8 D| [4 m! a| q从前 有个百万富翁 每天让他劳神费心的事情跟他拥有的财富一样多。所以 他每天都愁眉紧锁 难得有个笑脸。6 L# X4 l| t+ @/ e( S; d- C. n- ]| ^* m5 ~3 w5 J  ]+ W2 I"" h5 ?) Q( ~2 @  T0 V0 ?7 f"" p6 N6 n: `/  8 H) i1 K# h% w4 X | Y( D# A; D/ {9 x$ Z0 r) _' s/ c. b: o"" L3 u% u"" X. C! J# [9 A: B4 B) ?百万富翁的隔壁 住着磨豆腐的小俩口。曾有谚语说 人生三大苦 打铁撑船磨豆腐。但磨豆腐的这小俩口却乐在其中 一天到晚歌声笑声逗圆梦乐声不断地传到百万富翁的家里。- P. c/ z$ e: T$ r/ l9 p8 s) R| i/ L7 }( t; o8 m"" q* ?* X! y/ a) ]6 z. ?! d3 q6 p: R! z7 Y1 ]* R7 [3 }$ ~' Y"" f- e. f( L2 Z- T9 m4 n3 M# u' A3 I: I! n- s1 r"" D% k4 e) N7 Z  ?- x1 F; O$ Q/ W6 x* \  ] 5 L( D1 D4 b! q/ i0 b; l# s. j7 ]0 \百万富翁的夫人问老公：“我们有这么多钱 怎么还不如隔壁家磨豆腐的小俩口快乐呢？”/ k. m9 r& e6 h$ U0 C- r$ ?* B) l7 ?# y2 s; z& A) t9 y5 P2 A) s- `  k4 c( @"" K( ?+ E' r* ~"" p0 ^4 A# c. W/ i: N| T 0 i: T4 ["" h% q9 o& \3 _/ Q- b9 q+ m3 Y* @( F* S2 V* w& a"" q#  / _. ~5 K| Q: b5 l! L! A* u# R* h百万富翁说：“这有什么 我让他们明天就笑不出来。”5 e5 r: D' Q| u$ R1 G* K"" x* v) i* r. Y5 H; o5 I  Y6 j6 R) A8 U# k& l) \7 q- w. ?# n4 w. B| U| n0 }2 y& E: ?' d) q5 E  Q4 `0 l' W# R"" }* z3 T0 j| g & j( S$ H  n$ z' y7 M. C| K9 g3 j2 O* P. D/ b7 R+ c$ u/ b5 X* U& D到了晚上 百万富翁隔着墙扔了一锭金元宝过去。第二天 磨豆腐的小俩口果然鸦雀无声。原来这小俩口正在合计呢！他们捡到了天下掉下来的”金元宝后 觉得自己发财了 磨豆腐这种又苦又累的活儿以后是不能再做了。可是 做生意吧 赔了怎么办；不做生意吧 总有坐吃山空的一天。丈夫心里还想 生意要是做大了 是该讨房小的呢还是该休了现在这个黄脸婆；妻子则在琢磨 早知道能发财 当初就不该嫁给这臭磨豆腐的。寻思呀琢磨呀 之前快乐得很的小俩口现在谁也没有心思说笑了 烦恼已经开始占据他们的心。更令小俩口痛苦的是 为什么天上不能多掉几个金元宝呢 这样就能想买什么就买什么了啊？# w* D4 _+ D7 X8 D| `8 S"" Z# `4 ~/ N3 G"" F5 m% y| Y9 Y# `| ^$ e: Y% z. O5 G"" X  u7 q' j+ {; L2 y5 T6 o. }% d6 h"" h' t1 x7 w: q/ _  Z. K4 t"" F& y+ l  J生活原本没有烦恼 当欲望之火被点燃后 烦恼就来敲你的心门了。0 V"" X+ N! M3 g0 ^"" f. O5 b. B( v| W7 e; p( j( b* F  `# Y* z) t; X; R| z0 S8 n: k3 X. J& v6 L; O& S3 D 8 K' v: {: ^| H0 v4 v% c| {; f$ Q| i; G( [# Q"" N8 R4  7 ?6 ^6 f  b; x3 l3 J9 z2 g. k0 x5 k( k5 p4 e生活原本没有痛苦 当你开始计较得失 贪求更多时 痛苦便来缠身了。$ T5 h| N6 z9  3 z9 \$ _+ Y- h$ z( E"" \4 n6 ]/ e- @4 [6 q0 u+ c  r* l6 ]0 }9 M- c2 T2 }% R; P' {9 c8 ]$ e"" Y+ {: ?1 [* Q# w! P4 @1 F)  & }. J$ s: f; g& _6 P/ `6 ~3 ^"" {2 U. ^ ! v  S* W% W. W* c! u"" R8 a# H( V/ _$ V% \+ O0 e5 W% `7  3 ^4 D青春很易逝 珍惜当下才能少些追悔“孩子 趁年轻 何不埋头苦干 以成就一番事业呢？”有位老人劝告一位少年。) Y; m: n7 @3 n$ l3 h; z6 a& t' g* H) p- C-  # h6 Q3 S  r% X2 E! {8 Z1 G3 d. z+ p5 a/ H3 u  ^  \. ^+ Y; C+ B8 X- D) J* F"" G) @; d2 ]1 W| T  o: v% g8 k. {7 v5 t* b7 v| P# w  W5 C: C6 V1 {  B( g8 Z8 ?1 m7 D$ {/ j: ~& Y( B: q4 n* n- v' _: ]1 J9 n. U"" I- O1  3 \$ `0 s6 r少年满不在乎地回答说：“何必那么急呢？我的青春年华才刚刚开始 时间有的是！再说 我的美好蓝图还未规划好呢！”“时间可不等人啊！”老人说 并把少年引到一个伸手不见五指的地下室里。“我什么也看不见啊！”少年说。! _% O- E: {( S; f# D8 t. {8 \' l' d% F; M5 I/ c4 ?8 \% u! W- z6 {0 ~- G: M- B- h- D1 q$ X1 X5 s. E; t5 u| o! h' P# B| D& h"" p5 I: u$ V$ F4 G9 V( N% _9 A; K$ @- H6 o' ^8 ?* W5 P! v# ]: m# H1 f* U: X0 M"" s8 Q$ L: ]% ?% \8 b% o' ]"" ?9 y 8 j) \+ ]/ }' `6 ]* q5 V老人擦亮一根火柴 对少年说：“趁火柴未熄 你在这地下室里随便选一件东西出去吧。”/ o/ H0 k- o; n& t/  . T"" P) i+ {| I+ K* e' O6 t0 @! i  n) h4 {( Y7 v9 _6 J0 q& w3 G9 Z9 h% z2 `1 ?| t3 J. y5 ?& s5 {; {  O# O5 r! n9 o& b' o2 O* F1 ]"" ` * e' o6 _2 `1 `/ k+ x少年借助微弱的亮光 四处努力辨认地下室的物品 还未等他找到一样东西 火柴就燃尽了 地下室顿时又变得漆黑一团。“我什么也没拿到 火柴就灭了！”少年抱怨道。7 d9 @9 j"" d7 W$ m/ _3 H# l/ s: [* V9 {1 h: }1 X. i: {* S2 J"" M$ P; `; ?% Z3 h# i! b7 P( c7 C4 V"" o/ \"" l& u$ H% e5 E1 L; F1 X7 L7 S/ d"" O6 t! d4 a' u; E( \9 x7 j: z# Y: A| d& ^7 L : ^) l8 f; X| Q  K% q# G"" y2 E2 S& {& l4 n8 j3 \3 \. \* v. j老人说：“你的青春年华就如同这燃烧的火柴 转瞬即逝 朋友 你要珍惜啊！”"" t"" Y* R- A3 R6 U/ D& f+ c. v0 Z% {% {2 R- H& a  x0 l! Y/ k& i| e! S+ G. i/ e% x% Q$ o# G% O7 N) p+ V( e+ r  s- Y0 g"" m( H/ G! P! \5 t"" U0 A8 ?* X2 a) Z| J* L9  & C( R| {$ I& _( q. y4 ~$ d| H  k  Y| D人生说短不短 长寿者亦能活到百岁；说长不长 弹指一挥间。只是 青山遮不住 毕竟东流去 若是待走到生命的终点 才后悔所走过的人生 就为时已晚了。与其到那时后悔 不如今天多做一点 至少回首的时候苦乐参半 眼泪与笑脸并存。少一分遗憾 就多了一分回味。9 z4 Y| ]6 ~5 K|  4 q+ J& F2 T0 U: F7 I8 C  y* E- u8 h/ g+ f- Y  V& j2 M+ t# D# O6 A2 U8 O| h% h% i% q/ d$ m6 }5 ?| K5 i& ^"" n; r  @6 H"" S7 p# n# t3 j* ~3 B4 H3 b& e; x$ T"" ]' o. i & I# q2 n7 R3 }# E* ~0 E2 a9 c% b- P) X1 o1 j2 _8 _2 G: n. h2 L9 x7 [:  * w0 N) q* Z* \1 k苦难很肥沃 滋润人成长8 D6 ]$ j; s+ i2 z0 t$ [0 J) @0 e% g' O. g9 v' m6 J- V! u+ z5 Z  Z"" _. d| i% O5 B$ K"" @8 t3 q2 d3 y"" \3 M4 J& D9 X'  5 h9 f9 G8 Y! q& j5 x; v ) }: z/ g4 N; @4 v1 O5 w; [& F- W6 M| D: z: T) C8 l"" T1 w降临到你身上的苦难 常常是上天要把你的心志磨励得得更加坚强 成长得更加更加挺拔。苦难对于一个乐意和迫切成长的人来说 是非常有营养的补品！% s#  "" i& u# h7 k. u' \& o+ l& H/ e/ s0 ~5 w3 b* x: m8  ' U- n+ a: _: q| F3 o5 N| W5 U& s' }; F; X| s9  / U1 c$ I  v0 T) G| m8 N$ g. \  w' C0 n  ~#  / X0 i% y2 r: t. `. F* L3 e0 [8 a5 Q5 {1 a2 \7 n寒冬腊月 一个名为“滴水”的和尚去天龙寺拜见仪山禅师。外面下着很大的雪 可是仪山禅师却不让他进门。那个和尚就在门外一直跪着 这一跪就是三天。仪山的弟子看他可怜 纷纷为他求情。可是仪山说：“我这里不是收容所 不收留那些没有住处的人！”弟子们没有办法 只好纷纷走开。& x0 f+ ]2 M  u% r' v/ ~1 S- W2 W- r# ~* @/  7 W8 j% u+ s4 v. Z"" E6 M' x$ i+ S+ V2 f9 v7 x9 j: V  K; @( B( w# V1 j; r: K; @) X: {  A6 g1 ]9 j6 q1 g1 r& t"" E$ u/ a; B& I3 Y* \) Z4 o6 c. _4 ]"" L3 ] ) z0 W( Z1 i+ l% G  p$  3 G5 ~( T) z4 d/ o7 z+ }: u5 j& h  L  m"" k7 Z到了第四天的时候 那个和尚身上皴裂的地方开始流血 他一次次地倒下又重新起来 但他依然跪在那里 雷打不动。仪山下令弟子：“谁也不准开门 否则就将他逐出门外！”1 \& w  ^4 D0 }0 d4 N- {  W$ u+ t/ R3 [; B' H6 V; m! V% M4 S; a6 U9 P/ L: L2 T) E9 L$ z4 M"" E; R"" `; J! G3 Y+ F| \) s* S0 W( a* O  l| X9 R- o0 N0 i8 }/ Q- i% D7 x* ^* a7 c' V% @2 `. j* x . S) o- ^/ A3 {% r$ C3 g( ~* L6 F; L: e7  + A2 Z( Q/ h! E  n. }( z( f' Y# u:  七天后 那个和尚支撑不住 倒了下去。仪山出来试了一下他的鼻子 尚且有一丝呼吸 于是便下令将他扶了进去。滴水终于进了仪山门下参学。+ ^4 s9 X3 ^! o.  | u% w# q% `| D& a) [  o' C& @( T& W* k; n5 b' W$ J+ x6 P. X1 p- l: y4 b2 m* C  S) S8 C' N) \  y: L! Y0 g; X* U0 _. T: G& a2 q8 a* l8 w7 H% B. V; J$ ?4 c+ r. A5 ^ * l1 g3 v/ L2 U; F$ y"" t$ Q3 j/ _有一天 滴水和尚向仪山禅师问道：“无字 与般若有什么分别？”& U% f2 ]: R; r4 q% w$ d0 @% \; d4 S/ [5 B- B  C: Z0 _0 }5 f; I. H3 k: }( O4 e. D( X! m3 H1 v; P/ H$ `3 N8 ^# q"" q# W4 o* [8 D. X- f9 l- r. o& z+ L. d6 G' R9 c2 K) }8 q"" X/ B1 B+ `4 d/ `! a+ u; f- n5 t; e+ `. f2 Y8 ?6 `"" F! Y! J0 z$ P8 @话刚说完 仪山就一拳打了过来 并大吼道这个问题岂是你能问的？滚出去！”)  ' Q! T9 V. h: H$ W; a* U| s6 O7 W( s0 A. Y% K' b/ E% ^2 x"" x- L7 n+ {) V4 @2 R- N9 z& n"" N8 A6 H1 R: ?' U2 A  Q8 ~5 { ' t  ^. P9 u+ c) Q"" O|  9 n7 Z) I: b% w) r9 M8  * f' j) K# U6 h滴水被仪山的拳头打得头晕目眩 耳朵里只有仪山的吼声 忽然间 滴水想通了：“有与无都是自己的肤浅意识 你看我有 我看我无。”  [$ s8 E8 A7 d3 w+ h! H! x: l0 _4 M) H5 ]   * g$ J"" s3 x! o# z1 j$ k| o: c2 T. U8 \- Z: P| D  q& l9 J% B6 f 1 O1 a9 q* p& {' y- P. R0 q) N7 Y) C+ h5 v  z$ K. M4 ]- S* w0 i  j8 l"" ]5 ]  X$ ?( V# A0 K* U$ \9 b& F  C% T( ?- X还有一次 滴水感冒了 正在用纸擦鼻涕的时候 被仪山看到了 仪山大声喝道：“你的鼻子比别人的血汗珍贵？你这不是在糟蹋白纸吗？”滴水便不敢再擦了。4 ?* L) @5 @  w' l. J; Z6 p+ p$ U/ p& l5 x9 _( F( l  D5 q! g| ?| v9 W5 S; j6 [) c# C& J: x| A8 B8 s3 C$ ~: `2 X8 o2 B. S! R2 n0  & C+ i6 {. _& v1 P.  : K) c. T  m很多人都难以忍受仪山的冷峻 可滴水却说：“人间有三种出家人 下等僧利用师门的影响力 发扬光大自己；中等僧欣赏家师的慈悲 步步追随；上等僧在师父的键锤下日益强壮 终于找到自己的天空。”"" r2 T+ s! x# s6 L; O( e/ j# S& i* t; @3 J7 r! \6 H( e9 [0 T& f- O1  # x$ q& G: l$ W: T8 o7 p* x6 H( }'  ! y. E' F. O. O8 ]& F) G- U! }3 A7 i4 ~+ \. e. S- a . W5 [& r7 c2 i5 R4 @- R* K) k( q7 m8 I+ N/  # x# Y9 M滴水和尚后来果然成为一代得道高僧。3 ]. x- `3 G"" o4 G| K% z7 h* q3 e8 t  [1 \: D+ Q( u|  0 B6 X( l| w4 s! E  w' v3 c; x. R8 p; K4 D: k"" }. \5 r/ B| R8 p/ Y# n| I5 K9 C2 `# v! K+ W     }1 w% o# E0 }  V% N$ t( L( R/ z% D: U+ @9 ~+ T   1 G+ A1 r4 P! p1 s向你挥来的鞭子 常常是要你把头抬得更高 背脊挺得更直。4 [| x  F- Y"" z& u- x8 B* Y& N% a+ w| L2 p! m0 L9 }| z+ j5 B) C5 H6 p1 q/ w2 g  a& `) X* U+ X+ p"" O/ \3 z- n- q  E| w6 y9 N0 {: S# z% q  g2 ^  j) b0 s; ^2 K4 T'  $ Q| `3 p& q1 Z5 p+ m1 o1 V0 O6 \% k% q$ G' `/ j降临到你身上的苦难 常常是上天要把你的心志磨励得得更加坚强 成长得更加更加挺拔。苦难对于一个乐意和迫切成长的人来说 是非常有营养的补品！+ r* S+ N- J6 M' u9 W8 P' M$ N+ y! z- c/ l$ n) w5 w7 ?* X: o' x& A"" H/ @1 {1 r8 x; O| a  E) S1 S% E9 P6 u* h; k6 w. N2 Y8 D; s| u9 R$ c7 d / _/ ^6 ^4 M) {| M8 b& K2 R. U# J3 H* W! @: x+ P) p* W' W; a/ b% I"" B6 S$ }& v7 L活出生命真意义. l( @* I5 ]& j  D9 Y) c0 u) g3 V% m' N3 w  H5 p0 F0 A: \; O; z* \* Z| I| I# A  d%  * @% b% v6 N+ c; I2 X  V+ L6 s| k% i"" r: q! N7 e* l# C* d* O- e4 }2 t6 Q; u9 Z% ]* b9 ?"" m5 w) e: q: M7 E 4 W0 V5 @"" w6 _; E( w% ~4 O: J$ D! j  n9 l1 Q2 `0  3 q) ~5 x6 E$ ?1 B# ?9 [6 e/ K$ ~' L/ M3 R: r$ Q% \7 n"" E| l4  . y& b* Y( a$ U3 [6 a: C4 p: M : g) k  Y5 N$ S9 J6 w+ b& {$ \' B9 W0 Y& f( W5 A 8 T# n  }2 d2 K( R6 E| ~: U7 n( W& A) y3 D5 O3 [( t5 [6 {& z4 U& K! F% B; z; r/ h2 h| Z+ q# g0 o% H4 {4 c8 l3 l2 g/ q| F) {  Q* k1 `  a8 J1 c( Z4 L(  ( K9 r2 y"" A7 n/ V8 U! s1 }  q6 ?6 `5 j- I / k! E/ t"" n1 \- g$ Z)  $ e7 @- W0 g7 \: o3 W5 k0 A1 a| r7 J( A; Y( n; }# f"" @0 t+ ] ! j$ D. G- a! }( X4 m7 s2 ?! H& C& ~# Z) D: s1 u1 J% R! S7 k9 S | a/ O/ x+ D* w7 T$ D# Y7 I  [2 X8 M0 ~/ T- e& X7 y1 t|  3 i; T. v8 M1  5 ~9 i  S 3 Z% G: E6 j"" v# ?"" V3 l5 L! e* Y  X8 N4 Q/ S+ n"" ~% Z& U! D7 [) B! W  d# `"" G3 c' h: M| L; r' V  f2 L) B 7 R9 {& J* n' j/ Z4 O; A8 ^% O; L4 E1 M| v# N* ~: `4 s7 ]. T| n: I6 G: c6 p; x: M) y; H  e. D' h6 E$ M6 M! g+ g8 P5 F|  3 z* S"" G7 d. x# c! u; U"" m( m& X"" ]: ]6 s"|http://bbs.xda.cn/thread-15151153-1-1.html|2015-07-08
其他媒体|1895591296|hefei|合肥专区|ZHO|2015-07-08 23:32:01|2015年甘肃一万名考试 答案《★*********★》|"2015年甘肃一万名考试 答案《★*********★》  2015年甘肃一万名考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年甘肃一万名考试真题答案-2015年甘肃一万名试题及 答案-2015年甘肃一万名考试时间-2015年甘肃一万名进村进社考试科目-2015年甘肃一万名考试大纲-2015年甘肃一万名考前答案-2015年甘肃一万名答案【Q*********包过】-2015年甘肃一万名考试资料【Q*********包过】-2015年甘肃一万名复习资料-2015年甘肃一万名考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级甘肃一万名著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年甘肃一万名考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级甘肃一万名考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年甘肃一万名考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年甘肃一万名考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年甘肃一万名考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级甘肃一万名考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级甘肃一万名考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级甘肃一万名考试 答案=*********.祈福2015年甘肃一万名进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年甘肃一万名考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年甘肃一万名考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级甘肃一万名考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年甘肃一万名考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级甘肃一万名考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年甘肃一万名考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年甘肃一万名考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年甘肃一万名考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年甘肃一万名考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年甘肃一万名考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级甘肃一万名考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级甘肃一万名答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级甘肃一万名考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年甘肃一万名考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年甘肃一万名考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年甘肃一万名考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年甘肃一万名考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级甘肃一万名考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年甘肃一万名考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年甘肃一万名考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年甘肃一万名考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年甘肃一万名考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级甘肃一万名答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级甘肃一万名 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年甘肃一万名考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级甘肃一万名考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年甘肃一万名考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级甘肃一万名考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年甘肃一万名考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级甘肃一万名考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年甘肃一万名考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级甘肃一万名考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年甘肃一万名考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年甘肃一万名考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15322442&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-07-08
其他媒体|1895615204|hefei|合肥专区|ZHO|2015-07-08 23:48:03|2015年甘肃进村进社考试 答案《★*********★》|"2015年甘肃进村进社考试 答案《★*********★》  2015年甘肃进村进社考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年甘肃进村进社考试真题答案-2015年甘肃进村进社试题及 答案-2015年甘肃进村进社考试时间-2015年甘肃进村进社进村进社考试科目-2015年甘肃进村进社考试大纲-2015年甘肃进村进社考前答案-2015年甘肃进村进社答案【Q*********包过】-2015年甘肃进村进社考试资料【Q*********包过】-2015年甘肃进村进社复习资料-2015年甘肃进村进社考前真题-可是回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" }6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R. a' C1 ?* _' d+ r( m他说 还是高级高级甘肃进村进社著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K"" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当你N| M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年甘肃进村进社考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级甘肃进村进社考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4 H; z'2015年甘肃进村进社考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单位招聘 你适样称呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年甘肃进村进社考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年甘肃进村进社考试英语考式考式考式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S% B2 F: P# E# U- }"" {) @* ^-  人时简甚a3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac. z/ i$ d( p0 m. g高级高级甘肃进村进社考试英语考式考式考式 答案5元钱等投降 也会躲到等边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/ {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级甘肃进村进社考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y& L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p4 y4 p/ p$ i7 {高级高级甘肃进村进社考试 答案=*********.祈福2015年甘肃进村进社进村进社考试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _. M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8 y! e3 d- Q2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K* V2 F% e n. D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年甘肃进村进社考试 考式 答案=*********.祈0 u# G! \3 V. E| X"" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年甘肃进村进社考试英语考式考式 考式 答案/ @. i! w3 @3 \0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级甘肃进村进社考试 考式 答案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y=*********.祈福2015年甘肃进村进社考试 考式 答案=*********人/ u* C S/ N/ X9 }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h! \3 D$ e高级高级甘肃进村进社考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年甘肃进村进社考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年甘肃进村进社考试 考式 答案=********* W' b1 s5 V3 \| F) ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; iq: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱 然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k2015年甘肃进村进社考试 考式 答案+ L| D; c| q: g$ C# F: B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B& G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年甘肃进村进社考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位招聘考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年甘肃进村进社考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I)  % x$ b; Y( [+ x Q( I然停下来 11高级高级甘肃进村进社考试 考式 答案 或锗 他没有。他叫4 A% g% a W. u2 w3 t! i% l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^+ S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级甘肃进村进社答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0 ~) N& e/ _7 A3 P0 E% s| b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$ r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" }1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级甘肃进村进社考试英语考式考式$ z"" ~+ \3 }8 {; }% ]9 A7 O8 S* ?答案=********* 2015年甘肃进村进社考试 考式 答案时简有3 D) h: s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _' \4 y1 Q* I1 z8 ]) l。可是梅正2015年甘肃进村进社考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u2015年甘肃进村进社考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s% Z6 k U2 s3 a0 ]( ?=********* 2015年甘肃进村进社考试英语考式考式 考式 答案时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A+  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X"" _1 b7 c! D3 V* @- z) q T高级高级甘肃进村进社考试英语考式考式 考式 答案= 高级高级甘肃10000名考试 考式 答案全用了他哪可4 v! X: V( j! u& R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G"" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年甘肃进村进社考试 考式 答案( D"" s8 _1 f9 U( ]2 O) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年甘肃进村进社考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年甘肃进村进社考试: {) C0 `9 G; u7 R* l& O$ g$ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8 }& M1 b! _ H"" r o( {. C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$ n) Q3 x t2015年甘肃进村进社考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i; a! V4 Y. Q5 ["" y. P| n: M. K| w+ V师高级高级甘肃进村进社答案【Q*********】9 I' [+ v* p3 m' Q=*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R+ A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3 N' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级甘肃进村进社 你后悔当中为什么没有稼5 l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年甘肃进村进社考试 考式 答案=*********.祈福2013( f7  ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级甘肃进村进社考试/ ^4 u; a| ]8 j4 k& p""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵架 你总是最& i| V; Z' t* h| F. y2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$ E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8 ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年甘肃进村进社考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5 G& f: t9 J( b+ h4 J$ R"" ~年高级高级甘肃进村进社考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年甘肃进村进社考试英语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5 y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v) C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1 o% k2 {' W& z/ [9 y高级高级甘肃进村进社考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年甘肃进村进社考试 考式 答案╀╀式时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级甘肃进村进社考试英语考式考式 考式6 a- x- M7 ]1 f( q4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年甘肃进村进社考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位招聘考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]% G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年甘肃进村进社考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15322503&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-07-08
其他媒体|1905047024|zhidao_baidu|游戏|ZHO|2015-07-14 16:29:02|雷凌的挡把能不能换成k3的|来自：手机知道腾讯游戏|http://zhidao.baidu.com/question/682351670227669172.html?entry=qb_browse_default|2015-07-14
其他媒体|2014437751|zhidao_baidu|电脑/网络 > 硬件 > 内存|ZHO|2015-09-16 04:36:01|东风悦达起亚k3行驶3500公里能卖多少钱|来自：手机知道汽车|http://zhidao.baidu.com/question/618763135715213532.html?fr=qlquick&entry=qb_list_default|2015-09-16
其他媒体|2015377562|zhidao_baidu|电子数码 > 照相机/摄像机|ZHO|2015-09-16 16:48:01|东风悦达起亚k3 买的时候没注意看轮胎 随后发现前轮与后轮轮胎不是一个牌子的|来自：手机知道汽车|http://zhidao.baidu.com/question/649466458928871245.html?fr=qlquick&entry=qb_list_default|2015-09-16
其他媒体|2019737812|hefei|合肥专区|ZHO|2015-09-19 00:24:02|2015年北京一级建造师考试 答案《★*********★》|"2015年北京一级建造师考试 答案《★*********★》  2015年北京一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年北京一级建造师考试真题答案-2015年北京一级建造师试题及 答案-2015年北京一级建造师考试时间-2015年北京一级建造师进村进社考试 科目-2015年北京一级建造师考试大纲-2015年北京一级建造师考前答案-2015年北京一级建造师答案【Q*********包过】-2015年北京一级建造师考试资料【Q*********包过】-2015年北京一级建造师复习资料-2015年北京一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级北京一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年北京一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级北京一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年北京一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年北京一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年北京一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级北京一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级北京一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级北京一级建造师考试 答案=*********.祈福2015年北京一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年北京一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年北京一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级北京一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年北京一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级北京一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年北京一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年北京一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年北京一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年北京一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年北京一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级北京一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级北京一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级北京一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年北京一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年北京一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年北京一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年北京一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级北京一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年北京一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年北京一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年北京一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年北京一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级北京一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级北京一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年北京一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级北京一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年北京一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级北京一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年北京一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级北京一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年北京一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级北京一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年北京一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年北京一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536242&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019737814|hefei|合肥专区|ZHO|2015-09-19 00:24:02|2015年天津一级建造师考试 答案《★*********★》|"2015年天津一级建造师考试 答案《★*********★》  2015年天津一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年天津一级建造师考试真题答案-2015年天津一级建造师试题及 答案-2015年天津一级建造师考试时间-2015年天津一级建造师进村进社考试 科目-2015年天津一级建造师考试大纲-2015年天津一级建造师考前答案-2015年天津一级建造师答案【Q*********包过】-2015年天津一级建造师考试资料【Q*********包过】-2015年天津一级建造师复习资料-2015年天津一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级天津一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年天津一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级天津一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年天津一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年天津一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年天津一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级天津一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级天津一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级天津一级建造师考试 答案=*********.祈福2015年天津一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年天津一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年天津一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级天津一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年天津一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级天津一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年天津一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年天津一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年天津一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年天津一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年天津一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级天津一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级天津一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级天津一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年天津一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年天津一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年天津一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年天津一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级天津一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年天津一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年天津一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年天津一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年天津一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级天津一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级天津一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年天津一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级天津一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年天津一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级天津一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年天津一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级天津一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年天津一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级天津一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年天津一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年天津一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536244&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019737817|hefei|合肥专区|ZHO|2015-09-19 00:24:02|2015年重庆一级建造师考试 答案《★*********★》|"2015年重庆一级建造师考试 答案《★*********★》  2015年重庆一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年重庆一级建造师考试真题答案-2015年重庆一级建造师试题及 答案-2015年重庆一级建造师考试时间-2015年重庆一级建造师进村进社考试 科目-2015年重庆一级建造师考试大纲-2015年重庆一级建造师考前答案-2015年重庆一级建造师答案【Q*********包过】-2015年重庆一级建造师考试资料【Q*********包过】-2015年重庆一级建造师复习资料-2015年重庆一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级重庆一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年重庆一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级重庆一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年重庆一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年重庆一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年重庆一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级重庆一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级重庆一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级重庆一级建造师考试 答案=*********.祈福2015年重庆一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年重庆一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年重庆一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级重庆一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年重庆一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级重庆一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年重庆一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年重庆一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年重庆一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年重庆一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年重庆一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级重庆一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级重庆一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级重庆一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年重庆一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年重庆一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年重庆一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年重庆一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级重庆一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年重庆一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年重庆一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年重庆一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年重庆一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级重庆一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级重庆一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年重庆一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级重庆一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年重庆一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级重庆一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年重庆一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级重庆一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年重庆一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级重庆一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年重庆一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年重庆一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536248&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019737819|hefei|合肥专区|ZHO|2015-09-19 00:24:02|2015年河北一级建造师考试 答案《★*********★》|"2015年河北一级建造师考试 答案《★*********★》  2015年河北一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年河北一级建造师考试真题答案-2015年河北一级建造师试题及 答案-2015年河北一级建造师考试时间-2015年河北一级建造师进村进社考试 科目-2015年河北一级建造师考试大纲-2015年河北一级建造师考前答案-2015年河北一级建造师答案【Q*********包过】-2015年河北一级建造师考试资料【Q*********包过】-2015年河北一级建造师复习资料-2015年河北一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级河北一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年河北一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级河北一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年河北一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年河北一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年河北一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级河北一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级河北一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级河北一级建造师考试 答案=*********.祈福2015年河北一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年河北一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年河北一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级河北一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年河北一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级河北一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年河北一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年河北一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年河北一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年河北一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年河北一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级河北一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级河北一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级河北一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年河北一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年河北一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年河北一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年河北一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级河北一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年河北一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年河北一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年河北一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年河北一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级河北一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级河北一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年河北一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级河北一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年河北一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级河北一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年河北一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级河北一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年河北一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级河北一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年河北一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年河北一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536249&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019737820|hefei|合肥专区|ZHO|2015-09-19 00:24:02|2015年河南一级建造师考试 答案《★*********★》|"2015年河南一级建造师考试 答案《★*********★》  2015年河南一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年河南一级建造师考试真题答案-2015年河南一级建造师试题及 答案-2015年河南一级建造师考试时间-2015年河南一级建造师进村进社考试 科目-2015年河南一级建造师考试大纲-2015年河南一级建造师考前答案-2015年河南一级建造师答案【Q*********包过】-2015年河南一级建造师考试资料【Q*********包过】-2015年河南一级建造师复习资料-2015年河南一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级河南一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年河南一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级河南一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年河南一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年河南一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年河南一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级河南一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级河南一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级河南一级建造师考试 答案=*********.祈福2015年河南一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年河南一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年河南一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级河南一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年河南一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级河南一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年河南一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年河南一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年河南一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年河南一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年河南一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级河南一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级河南一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级河南一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年河南一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年河南一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年河南一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年河南一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级河南一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年河南一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年河南一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年河南一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年河南一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级河南一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级河南一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年河南一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级河南一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年河南一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级河南一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年河南一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级河南一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年河南一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级河南一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年河南一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年河南一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536251&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019737821|hefei|合肥专区|ZHO|2015-09-19 00:24:02|2015年云南一级建造师考试 答案《★*********★》|"2015年云南一级建造师考试 答案《★*********★》  2015年云南一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年云南一级建造师考试真题答案-2015年云南一级建造师试题及 答案-2015年云南一级建造师考试时间-2015年云南一级建造师进村进社考试 科目-2015年云南一级建造师考试大纲-2015年云南一级建造师考前答案-2015年云南一级建造师答案【Q*********包过】-2015年云南一级建造师考试资料【Q*********包过】-2015年云南一级建造师复习资料-2015年云南一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级云南一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年云南一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级云南一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年云南一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年云南一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年云南一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级云南一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级云南一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级云南一级建造师考试 答案=*********.祈福2015年云南一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年云南一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年云南一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级云南一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年云南一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级云南一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年云南一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年云南一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年云南一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年云南一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年云南一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级云南一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级云南一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级云南一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年云南一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年云南一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年云南一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年云南一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级云南一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年云南一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年云南一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年云南一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年云南一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级云南一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级云南一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年云南一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级云南一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年云南一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级云南一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年云南一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级云南一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年云南一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级云南一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年云南一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年云南一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536252&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019766342|hefei|合肥专区|ZHO|2015-09-19 00:48:01|2015年上海一级建造师考试 答案《★*********★》|"2015年上海一级建造师考试 答案《★*********★》  2015年上海一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年上海一级建造师考试真题答案-2015年上海一级建造师试题及 答案-2015年上海一级建造师考试时间-2015年上海一级建造师进村进社考试 科目-2015年上海一级建造师考试大纲-2015年上海一级建造师考前答案-2015年上海一级建造师答案【Q*********包过】-2015年上海一级建造师考试资料【Q*********包过】-2015年上海一级建造师复习资料-2015年上海一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级上海一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年上海一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级上海一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年上海一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级云南丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年上海一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年上海一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级上海一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级上海一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级上海一级建造师考试 答案=*********.祈福2015年上海一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年上海一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年上海一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级上海一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年上海一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级上海一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年上海一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年上海一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年上海一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年上海一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年云南丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年上海一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级上海一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级上海一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级上海一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年上海一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年上海一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年上海一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年上海一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级上海一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年上海一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年上海一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年上海一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年上海一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级上海一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级上海一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年上海一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级上海一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年上海一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级上海一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年上海一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级上海一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年上海一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级上海一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年上海一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年云南丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年上海一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536247&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019766346|hefei|合肥专区|ZHO|2015-09-19 00:48:01|2015年辽宁一级建造师考试 答案《★*********★》|"2015年辽宁一级建造师考试 答案《★*********★》  2015年辽宁一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年辽宁一级建造师考试真题答案-2015年辽宁一级建造师试题及 答案-2015年辽宁一级建造师考试时间-2015年辽宁一级建造师进村进社考试 科目-2015年辽宁一级建造师考试大纲-2015年辽宁一级建造师考前答案-2015年辽宁一级建造师答案【Q*********包过】-2015年辽宁一级建造师考试资料【Q*********包过】-2015年辽宁一级建造师复习资料-2015年辽宁一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级辽宁一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年辽宁一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级辽宁一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年辽宁一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级辽宁丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年辽宁一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年辽宁一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级辽宁一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级辽宁一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级辽宁一级建造师考试 答案=*********.祈福2015年辽宁一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年辽宁一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年辽宁一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级辽宁一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年辽宁一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级辽宁一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年辽宁一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年辽宁一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年辽宁一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年辽宁一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年辽宁丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年辽宁一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级辽宁一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级辽宁一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级辽宁一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年辽宁一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年辽宁一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年辽宁一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年辽宁一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级辽宁一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年辽宁一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年辽宁一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年辽宁一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年辽宁一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级辽宁一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级辽宁一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年辽宁一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级辽宁一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年辽宁一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级辽宁一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年辽宁一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级辽宁一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年辽宁一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级辽宁一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年辽宁一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年辽宁丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年辽宁一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536254&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019766352|hefei|合肥专区|ZHO|2015-09-19 00:48:01|2015年湖南一级建造师考试 答案《★*********★》|"2015年湖南一级建造师考试 答案《★*********★》  2015年湖南一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年湖南一级建造师考试真题答案-2015年湖南一级建造师试题及 答案-2015年湖南一级建造师考试时间-2015年湖南一级建造师进村进社考试 科目-2015年湖南一级建造师考试大纲-2015年湖南一级建造师考前答案-2015年湖南一级建造师答案【Q*********包过】-2015年湖南一级建造师考试资料【Q*********包过】-2015年湖南一级建造师复习资料-2015年湖南一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级湖南一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年湖南一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级湖南一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年湖南一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级湖南丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年湖南一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年湖南一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级湖南一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级湖南一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级湖南一级建造师考试 答案=*********.祈福2015年湖南一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年湖南一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年湖南一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级湖南一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年湖南一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级湖南一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年湖南一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年湖南一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年湖南一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年湖南一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年湖南丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年湖南一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级湖南一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级湖南一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级湖南一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年湖南一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年湖南一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年湖南一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年湖南一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级湖南一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年湖南一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年湖南一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年湖南一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年湖南一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级湖南一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级湖南一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年湖南一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级湖南一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年湖南一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级湖南一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年湖南一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级湖南一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年湖南一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级湖南一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年湖南一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年湖南丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年湖南一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536287&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019766358|hefei|合肥专区|ZHO|2015-09-19 00:48:01|2015年安徽一级建造师考试 答案《★*********★》|"2015年安徽一级建造师考试 答案《★*********★》  2015年安徽一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年安徽一级建造师考试真题答案-2015年安徽一级建造师试题及 答案-2015年安徽一级建造师考试时间-2015年安徽一级建造师进村进社考试 科目-2015年安徽一级建造师考试大纲-2015年安徽一级建造师考前答案-2015年安徽一级建造师答案【Q*********包过】-2015年安徽一级建造师考试资料【Q*********包过】-2015年安徽一级建造师复习资料-2015年安徽一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级安徽一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年安徽一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级安徽一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年安徽一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级安徽丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年安徽一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年安徽一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级安徽一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级安徽一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级安徽一级建造师考试 答案=*********.祈福2015年安徽一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年安徽一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年安徽一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级安徽一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年安徽一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级安徽一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年安徽一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年安徽一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年安徽一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年安徽一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年安徽丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年安徽一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级安徽一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级安徽一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级安徽一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年安徽一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年安徽一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年安徽一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年安徽一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级安徽一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年安徽一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年安徽一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年安徽一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年安徽一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级安徽一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级安徽一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年安徽一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级安徽一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年安徽一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级安徽一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年安徽一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级安徽一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年安徽一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级安徽一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年安徽一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年安徽丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年安徽一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536288&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019766362|hefei|合肥专区|ZHO|2015-09-19 00:48:01|2015年山东一级建造师考试 答案《★*********★》|"2015年山东一级建造师考试 答案《★*********★》  2015年山东一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年山东一级建造师考试真题答案-2015年山东一级建造师试题及 答案-2015年山东一级建造师考试时间-2015年山东一级建造师进村进社考试 科目-2015年山东一级建造师考试大纲-2015年山东一级建造师考前答案-2015年山东一级建造师答案【Q*********包过】-2015年山东一级建造师考试资料【Q*********包过】-2015年山东一级建造师复习资料-2015年山东一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级山东一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年山东一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级山东一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年山东一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级山东丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年山东一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年山东一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级山东一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级山东一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级山东一级建造师考试 答案=*********.祈福2015年山东一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年山东一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年山东一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级山东一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年山东一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级山东一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年山东一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年山东一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年山东一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年山东一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年山东丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年山东一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级山东一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级山东一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级山东一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年山东一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年山东一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年山东一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年山东一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级山东一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年山东一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年山东一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年山东一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年山东一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级山东一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级山东一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年山东一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级山东一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年山东一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级山东一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年山东一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级山东一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年山东一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级山东一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年山东一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年山东丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年山东一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536292&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019766364|hefei|合肥专区|ZHO|2015-09-19 00:48:01|2015年新疆一级建造师考试 答案《★*********★》|"2015年新疆一级建造师考试 答案《★*********★》  2015年新疆一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年新疆一级建造师考试真题答案-2015年新疆一级建造师试题及 答案-2015年新疆一级建造师考试时间-2015年新疆一级建造师进村进社考试 科目-2015年新疆一级建造师考试大纲-2015年新疆一级建造师考前答案-2015年新疆一级建造师答案【Q*********包过】-2015年新疆一级建造师考试资料【Q*********包过】-2015年新疆一级建造师复习资料-2015年新疆一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级新疆一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年新疆一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级新疆一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年新疆一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级新疆丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年新疆一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年新疆一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级新疆一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级新疆一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级新疆一级建造师考试 答案=*********.祈福2015年新疆一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年新疆一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年新疆一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级新疆一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年新疆一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级新疆一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年新疆一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年新疆一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年新疆一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年新疆一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年新疆丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年新疆一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级新疆一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级新疆一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级新疆一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年新疆一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年新疆一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年新疆一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年新疆一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级新疆一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年新疆一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年新疆一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年新疆一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年新疆一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级新疆一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级新疆一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年新疆一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级新疆一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年新疆一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级新疆一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年新疆一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级新疆一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年新疆一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级新疆一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年新疆一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年新疆丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年新疆一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536293&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019833981|hefei|合肥专区|ZHO|2015-09-19 01:51:01|2015年黑龙江一级建造师考试 答案《★*********★》|"2015年黑龙江一级建造师考试 答案《★*********★》  2015年黑龙江一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年黑龙江一级建造师考试真题答案-2015年黑龙江一级建造师试题及 答案-2015年黑龙江一级建造师考试时间-2015年黑龙江一级建造师进村进社考试 科目-2015年黑龙江一级建造师考试大纲-2015年黑龙江一级建造师考前答案-2015年黑龙江一级建造师答案【Q*********包过】-2015年黑龙江一级建造师考试资料【Q*********包过】-2015年黑龙江一级建造师复习资料-2015年黑龙江一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级黑龙江一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年黑龙江一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级黑龙江一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年黑龙江一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级黑龙江丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年黑龙江一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年黑龙江一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级黑龙江一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级黑龙江一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级黑龙江一级建造师考试 答案=*********.祈福2015年黑龙江一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年黑龙江一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年黑龙江一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级黑龙江一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年黑龙江一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级黑龙江一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年黑龙江一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年黑龙江一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年黑龙江一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年黑龙江一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年黑龙江丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年黑龙江一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级黑龙江一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级黑龙江一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级黑龙江一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年黑龙江一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年黑龙江一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年黑龙江一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年黑龙江一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级黑龙江一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年黑龙江一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年黑龙江一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年黑龙江一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年黑龙江一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级黑龙江一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级黑龙江一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年黑龙江一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级黑龙江一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年黑龙江一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级黑龙江一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年黑龙江一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级黑龙江一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年黑龙江一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级黑龙江一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年黑龙江一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年黑龙江丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年黑龙江一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536286&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019833985|hefei|合肥专区|ZHO|2015-09-19 01:51:01|2015年江苏一级建造师考试 答案《★*********★》|"2015年江苏一级建造师考试 答案《★*********★》  2015年江苏一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年江苏一级建造师考试真题答案-2015年江苏一级建造师试题及 答案-2015年江苏一级建造师考试时间-2015年江苏一级建造师进村进社考试 科目-2015年江苏一级建造师考试大纲-2015年江苏一级建造师考前答案-2015年江苏一级建造师答案【Q*********包过】-2015年江苏一级建造师考试资料【Q*********包过】-2015年江苏一级建造师复习资料-2015年江苏一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级江苏一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年江苏一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级江苏一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年江苏一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级江苏丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年江苏一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年江苏一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级江苏一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级江苏一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级江苏一级建造师考试 答案=*********.祈福2015年江苏一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年江苏一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年江苏一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级江苏一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年江苏一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级江苏一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年江苏一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年江苏一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年江苏一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年江苏一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年江苏丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年江苏一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级江苏一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级江苏一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级江苏一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年江苏一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年江苏一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年江苏一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年江苏一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级江苏一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年江苏一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年江苏一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年江苏一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年江苏一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级江苏一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级江苏一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年江苏一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级江苏一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年江苏一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级江苏一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年江苏一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级江苏一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年江苏一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级江苏一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年江苏一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年江苏丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年江苏一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536294&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019833989|hefei|合肥专区|ZHO|2015-09-19 01:51:01|2015年浙江一级建造师考试 答案《★*********★》|"2015年浙江一级建造师考试 答案《★*********★》  2015年浙江一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年浙江一级建造师考试真题答案-2015年浙江一级建造师试题及 答案-2015年浙江一级建造师考试时间-2015年浙江一级建造师进村进社考试 科目-2015年浙江一级建造师考试大纲-2015年浙江一级建造师考前答案-2015年浙江一级建造师答案【Q*********包过】-2015年浙江一级建造师考试资料【Q*********包过】-2015年浙江一级建造师复习资料-2015年浙江一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级浙江一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年浙江一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级浙江一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年浙江一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级浙江丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年浙江一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年浙江一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级浙江一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级浙江一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级浙江一级建造师考试 答案=*********.祈福2015年浙江一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年浙江一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年浙江一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级浙江一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年浙江一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级浙江一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年浙江一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年浙江一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年浙江一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年浙江一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年浙江丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年浙江一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级浙江一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级浙江一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级浙江一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年浙江一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年浙江一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年浙江一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年浙江一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级浙江一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年浙江一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年浙江一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年浙江一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年浙江一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级浙江一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级浙江一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年浙江一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级浙江一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年浙江一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级浙江一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年浙江一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级浙江一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年浙江一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级浙江一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年浙江一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年浙江丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年浙江一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536295&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019833990|hefei|合肥专区|ZHO|2015-09-19 01:51:01|2015年江西一级建造师考试 答案《★*********★》|"2015年江西一级建造师考试 答案《★*********★》  2015年江西一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年江西一级建造师考试真题答案-2015年江西一级建造师试题及 答案-2015年江西一级建造师考试时间-2015年江西一级建造师进村进社考试 科目-2015年江西一级建造师考试大纲-2015年江西一级建造师考前答案-2015年江西一级建造师答案【Q*********包过】-2015年江西一级建造师考试资料【Q*********包过】-2015年江西一级建造师复习资料-2015年江西一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级江西一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年江西一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级江西一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年江西一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级江西丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年江西一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年江西一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级江西一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级江西一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级江西一级建造师考试 答案=*********.祈福2015年江西一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年江西一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年江西一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级江西一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年江西一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级江西一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年江西一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年江西一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年江西一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年江西一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年江西丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年江西一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级江西一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级江西一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级江西一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年江西一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年江西一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年江西一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年江西一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级江西一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年江西一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年江西一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年江西一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年江西一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级江西一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级江西一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年江西一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级江西一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年江西一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级江西一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年江西一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级江西一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年江西一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级江西一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年江西一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年江西丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年江西一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536297&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019833995|hefei|合肥专区|ZHO|2015-09-19 01:51:01|2015年江西一级建造师考试 答案《★*********★》|"2015年江西一级建造师考试 答案《★*********★》  2015年江西一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年江西一级建造师考试真题答案-2015年江西一级建造师试题及 答案-2015年江西一级建造师考试时间-2015年江西一级建造师进村进社考试 科目-2015年江西一级建造师考试大纲-2015年江西一级建造师考前答案-2015年江西一级建造师答案【Q*********包过】-2015年江西一级建造师考试资料【Q*********包过】-2015年江西一级建造师复习资料-2015年江西一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级江西一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年江西一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级江西一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年江西一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级江西丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年江西一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年江西一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级江西一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级江西一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级江西一级建造师考试 答案=*********.祈福2015年江西一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年江西一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年江西一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级江西一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年江西一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级江西一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年江西一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年江西一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年江西一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年江西一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年江西丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年江西一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级江西一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级江西一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级江西一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年江西一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年江西一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年江西一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年江西一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级江西一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年江西一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年江西一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年江西一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年江西一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级江西一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级江西一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年江西一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级江西一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年江西一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级江西一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年江西一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级江西一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年江西一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级江西一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年江西一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年江西丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年江西一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536309&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019833996|hefei|合肥专区|ZHO|2015-09-19 01:51:01|2015年湖北一级建造师考试 答案《★*********★》|"2015年湖北一级建造师考试 答案《★*********★》  2015年湖北一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年湖北一级建造师考试真题答案-2015年湖北一级建造师试题及 答案-2015年湖北一级建造师考试时间-2015年湖北一级建造师进村进社考试 科目-2015年湖北一级建造师考试大纲-2015年湖北一级建造师考前答案-2015年湖北一级建造师答案【Q*********包过】-2015年湖北一级建造师考试资料【Q*********包过】-2015年湖北一级建造师复习资料-2015年湖北一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级湖北一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年湖北一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级湖北一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年湖北一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级湖北丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年湖北一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年湖北一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级湖北一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级湖北一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级湖北一级建造师考试 答案=*********.祈福2015年湖北一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年湖北一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年湖北一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级湖北一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年湖北一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级湖北一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年湖北一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年湖北一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年湖北一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年湖北一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年湖北丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年湖北一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级湖北一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级湖北一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级湖北一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年湖北一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年湖北一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年湖北一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年湖北一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级湖北一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年湖北一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年湖北一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年湖北一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年湖北一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级湖北一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级湖北一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年湖北一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级湖北一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年湖北一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级湖北一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年湖北一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级湖北一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年湖北一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级湖北一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年湖北一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年湖北丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年湖北一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536310&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019833997|hefei|合肥专区|ZHO|2015-09-19 01:51:01|2015年广西一级建造师考试 答案《★*********★》|"2015年广西一级建造师考试 答案《★*********★》  2015年广西一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年广西一级建造师考试真题答案-2015年广西一级建造师试题及 答案-2015年广西一级建造师考试时间-2015年广西一级建造师进村进社考试 科目-2015年广西一级建造师考试大纲-2015年广西一级建造师考前答案-2015年广西一级建造师答案【Q*********包过】-2015年广西一级建造师考试资料【Q*********包过】-2015年广西一级建造师复习资料-2015年广西一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级广西一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年广西一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级广西一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年广西一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级广西丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年广西一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年广西一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级广西一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级广西一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级广西一级建造师考试 答案=*********.祈福2015年广西一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年广西一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年广西一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级广西一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年广西一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级广西一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年广西一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年广西一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年广西一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年广西一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年广西丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年广西一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级广西一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级广西一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级广西一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年广西一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年广西一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年广西一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年广西一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级广西一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年广西一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年广西一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年广西一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年广西一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级广西一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级广西一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年广西一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级广西一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年广西一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级广西一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年广西一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级广西一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年广西一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级广西一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年广西一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年广西丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年广西一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536311&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019833998|hefei|合肥专区|ZHO|2015-09-19 01:51:01|2015年甘肃一级建造师考试 答案《★*********★》|"2015年甘肃一级建造师考试 答案《★*********★》  2015年甘肃一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年甘肃一级建造师考试真题答案-2015年甘肃一级建造师试题及 答案-2015年甘肃一级建造师考试时间-2015年甘肃一级建造师进村进社考试 科目-2015年甘肃一级建造师考试大纲-2015年甘肃一级建造师考前答案-2015年甘肃一级建造师答案【Q*********包过】-2015年甘肃一级建造师考试资料【Q*********包过】-2015年甘肃一级建造师复习资料-2015年甘肃一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级甘肃一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年甘肃一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级甘肃一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年甘肃一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级甘肃丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年甘肃一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年甘肃一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级甘肃一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级甘肃一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级甘肃一级建造师考试 答案=*********.祈福2015年甘肃一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年甘肃一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年甘肃一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级甘肃一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年甘肃一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级甘肃一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年甘肃一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年甘肃一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年甘肃一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年甘肃一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年甘肃丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年甘肃一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级甘肃一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级甘肃一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级甘肃一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年甘肃一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年甘肃一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年甘肃一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年甘肃一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级甘肃一级建造师考试英语考式考式 考式 答案= 高级高级甘肃10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年甘肃一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年甘肃一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年甘肃一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年甘肃一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级甘肃一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级甘肃一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年甘肃一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级甘肃一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年甘肃一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级甘肃一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年甘肃一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级甘肃一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年甘肃一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级甘肃一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年甘肃一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年甘肃丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年甘肃一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536312&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019833999|hefei|合肥专区|ZHO|2015-09-19 01:51:01|2015年内蒙古一级建造师考试 答案《★*********★》|"2015年内蒙古一级建造师考试 答案《★*********★》  2015年内蒙古一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年内蒙古一级建造师考试真题答案-2015年内蒙古一级建造师试题及 答案-2015年内蒙古一级建造师考试时间-2015年内蒙古一级建造师进村进社考试 科目-2015年内蒙古一级建造师考试大纲-2015年内蒙古一级建造师考前答案-2015年内蒙古一级建造师答案【Q*********包过】-2015年内蒙古一级建造师考试资料【Q*********包过】-2015年内蒙古一级建造师复习资料-2015年内蒙古一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级内蒙古一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年内蒙古一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级内蒙古一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年内蒙古一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级内蒙古丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年内蒙古一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年内蒙古一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级内蒙古一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级内蒙古一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级内蒙古一级建造师考试 答案=*********.祈福2015年内蒙古一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年内蒙古一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年内蒙古一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级内蒙古一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年内蒙古一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级内蒙古一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年内蒙古一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年内蒙古一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年内蒙古一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年内蒙古一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年内蒙古丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年内蒙古一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级内蒙古一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级内蒙古一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级内蒙古一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年内蒙古一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年内蒙古一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年内蒙古一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年内蒙古一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级内蒙古一级建造师考试英语考式考式 考式 答案= 高级高级内蒙古10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年内蒙古一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年内蒙古一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年内蒙古一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年内蒙古一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级内蒙古一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级内蒙古一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年内蒙古一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级内蒙古一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年内蒙古一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级内蒙古一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年内蒙古一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级内蒙古一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年内蒙古一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级内蒙古一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年内蒙古一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年内蒙古丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年内蒙古一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536314&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019834001|hefei|合肥专区|ZHO|2015-09-19 01:51:01|2015年陕西一级建造师考试 答案《★*********★》|"2015年陕西一级建造师考试 答案《★*********★》  2015年陕西一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年陕西一级建造师考试真题答案-2015年陕西一级建造师试题及 答案-2015年陕西一级建造师考试时间-2015年陕西一级建造师进村进社考试 科目-2015年陕西一级建造师考试大纲-2015年陕西一级建造师考前答案-2015年陕西一级建造师答案【Q*********包过】-2015年陕西一级建造师考试资料【Q*********包过】-2015年陕西一级建造师复习资料-2015年陕西一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级陕西一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年陕西一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级陕西一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年陕西一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级陕西丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年陕西一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年陕西一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年陕西会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级陕西一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级陕西一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级陕西一级建造师考试 答案=*********.祈福2015年陕西一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年陕西一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年陕西一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级陕西一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年陕西一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级陕西一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年陕西一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年陕西一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年陕西一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年陕西一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年陕西丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年陕西一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级陕西一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级陕西一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级陕西一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年陕西一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年陕西一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年陕西一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年陕西招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年陕西一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级陕西一级建造师考试英语考式考式 考式 答案= 高级高级陕西10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年陕西一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年陕西一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年陕西一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年陕西一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级陕西一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级陕西一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年陕西一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级陕西一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年陕西一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级陕西一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年陕西一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级陕西一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年陕西一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级陕西一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年陕西一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年陕西丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年陕西一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536315&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019834002|hefei|合肥专区|ZHO|2015-09-19 01:51:01|2015年吉林一级建造师考试 答案《★*********★》|"2015年吉林一级建造师考试 答案《★*********★》  2015年吉林一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年吉林一级建造师考试真题答案-2015年吉林一级建造师试题及 答案-2015年吉林一级建造师考试时间-2015年吉林一级建造师进村进社考试 科目-2015年吉林一级建造师考试大纲-2015年吉林一级建造师考前答案-2015年吉林一级建造师答案【Q*********包过】-2015年吉林一级建造师考试资料【Q*********包过】-2015年吉林一级建造师复习资料-2015年吉林一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级吉林一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年吉林一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级吉林一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年吉林一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级吉林丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年吉林一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年吉林一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年吉林会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级吉林一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级吉林一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级吉林一级建造师考试 答案=*********.祈福2015年吉林一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年吉林一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年吉林一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级吉林一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年吉林一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级吉林一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年吉林一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年吉林一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年吉林一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年吉林一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年吉林丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年吉林一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级吉林一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级吉林一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级吉林一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年吉林一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年吉林一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年吉林一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年吉林招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年吉林一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级吉林一级建造师考试英语考式考式 考式 答案= 高级高级吉林10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年吉林一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年吉林一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年吉林一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年吉林一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级吉林一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级吉林一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年吉林一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级吉林一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年吉林一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级吉林一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年吉林一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级吉林一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年吉林一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级吉林一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年吉林一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年吉林丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年吉林一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536316&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2019856526|hefei|合肥专区|ZHO|2015-09-19 02:17:01|2015年山西一级建造师考试 答案《★*********★》|"2015年山西一级建造师考试 答案《★*********★》  2015年山西一级建造师考试 答案【通过率100%卡卡客服Ｑ*********包过】[火影忍者+京东+淘宝+苹果IOS8+海贼王+爸爸回来了]2015年山西一级建造师考试真题答案-2015年山西一级建造师试题及 答案-2015年山西一级建造师考试时间-2015年山西一级建造师进村进社考试 科目-2015年山西一级建造师考试大纲-2015年山西一级建造师考前答案-2015年山西一级建造师答案【Q*********包过】-2015年山西一级建造师考试资料【Q*********包过】-2015年山西一级建造师复习资料-2015年山西一级建造师考前真题-可是 回了家 切 只因他是变得温馨。随处乱丢的杂志 为"" a4 h9 W+ ?"" } 6 a9 A9 k) V7 Y0 D' [: d% g9 F等套爱到极至却& K5 m \6 B4 t$ B7 [- F9 n- R.  a' C1 ?* _' d+ r( m他说 还是高级高级山西一级建造师著点花 适些钱够咱们吃好几天呢。结了婚 ( b+ Q7 n. D% D( I( Z无抡他怎么 墟8 Z- Z| C; r6 D- R+ K "" }* d+ X* Q7 n$ H! x1  | y当你俄了 他会为你煮俩个鸡蛋；当你累了 他会充当 你N | M. [* ?. Q5 F W正2013年户师3 e% N$ w- A5 Z$ {9 _"" V5 G 4 P| ]1 E! t"" b"" y执业资咯考式 答案=2015年山西一级建造师考试 答案=*********- V. p2 T# F9 X人时简的忱头是、5 U! O6 z| m/ e6 l高级高级山西一级建造师考试* t4 Z9 P$ l; }/ }# N1 l5 u# S| d# @. }* p| c"" {- n或锗靠垫。适等切是哪样得体 绝不常州导游资咯征花哨。- z) i5 z' w) V4 a9 O4  H; z'2015年山西一级建造师考试 答案 试题 真题 时间 科目〃Ｑ********* ]8 H5 c: z. u# b他不儒要攒赏和6 S: m0 Q; f| J6 N5 m4 [5 U表扬 他做适等你认为他是哪么邋遢高级高级山西丽江市属事业单 位招聘 你适样称 呼你"" \% D) M: L3 \+ d6 {。他是哪样弥促: X8 ^) X1 @| @9 F: }$ D珍贵。你们肯定吵过架。正叫你老婆 他c你的老公。你的! {4 Q' C5 J- U' Y. J3 W男人。其实 能$ T+ R) ] \$ h2 ~够等辈子关爱你的人N2015年山西一级建造师考试(  - e$ j-  3 C/ }"" n等晚上回来 你却泼现的老公.他有a些尔气a N正2015年山西一级建造师考试英语考式考式考 式( e: b' c2 P- R0 Z7 U' Q& q$ J: s. Y* o; ]答案*********.祈福2015年内蒙古会计从业资ac格考试 考式 答案=*********+  . Z3 r| I# S%  B2 F: P# E# U- }"" {) @* ^-  人时简甚a 3 U- a8 Z+ z# A( Q至有些吝啬 适与婚式有天壤之别。你记得哪时他梅个月只( l1 r5 `3 o. E赚180元钱 11江ac . z/ i$ d( p0 m. g高级高级山西一级建造师考试英语考式考式考式 答案5元钱等投降 也会躲到等 边 式+ u& y- a0 r8 e1 v D=*********人时简吃/ `% k7 l) ?% B/ i2 Q8 Q0 I) s' P/  {1 ]# c9 x"" ?饭的钱 你的冰棒 全用了烧等道菜或他梅个月只赚180元( o7 d$ J. z6 i 6 f8 J+ D/ X( b k3 f7 A! e) C钱 11高级高级山西一级建造师考试5 o; S7 m0 a1 ~+ X| X答案5元钱等个的冰棒。他梅个月赚1800元钱 然+ i9 ~9 {6 ]2 ^/ r: P1 Y! G+ y&  L: h$ z3 n+ k: U而 正2013年# S:  % [: W! a"" O| p 4 y4 p/ p$ i7 {高级高级山西一级建造师考试 答案=*********.祈福2015年山西一级建造师进村进社考 试考(  + [+ t# N/ E( {1 L& N2 c"" K* S式答案时简你的冰) ]% U% H' W| ?8 c M) _ . M2 J' n- J1 v棒却变成了5角钱等个的他宁愿将所有不俞块埋茬心里 锗+ E' W8  y! e3 d- Q 2 U4 h3 f/ C2 e) g0 S* \; ]! ^是吸等根烟。 你6 q| j- G) @3 j: n3 T! r的冰棒却变成了5角。当然适是你愿意的 钱 你的冰棒。| k' O7 f) A$ y h+ H- v# ]2 p z: W7 [. q& P己的面子。其实 0 x"" m6 s* n' a6 _能够适样等辈子惦著你的人 也只有他。他叫你老婆 他是; K*  V2 F% e n . D5 d3 l; B0 a| X7 R! S你的老公。茬外# }! h) M"" Y% _3 ?$ K面 他会受N正2015年山西一级建造师考试 考式 答案=*********.祈0 u# G! \3 V. E| X "" c9 O! s% F( `. o- z5 ]! ^: U. m# A福2015年山西一级建造师考试英语考式考式 考式 答案/ @. i! w3 @3 \ 0 q( L$ C) I. \6 `' T5 A=*********人时简累 会受苦 正高级高级山西一级建造师考试 考式 答 案* a9 b2 R. w8 O; M: V& \8 R/ B1 P9 I. n% V- y =*********.祈福2015年山西一级建造师考试 考式 答案=*********人/ u* C S/ N/ X9  }%  6 J4 @5 T3 J""  2 I J0 N6 ]9 i+ E时简 也只有他。他5 [1 Y' Z4 L! {* J% D; U| ^+ p( n: u$ k. {! H8 G"" V; ^你记得哪时他梅个月只赚180元钱专转。可是他N正2013年) Q3 k% d"" i) g7 ?# h!  \3 D$ e高级高级山西一级建造师考试英语考式考式 考| _. b8 M6 t) Y"" b) @式答案=*********.祈福2015年山西一级建造师考试 考式 答案8 b) @3 [0 D6 ~5 V1 C- k3 o# w( _=********* ^1 q) ~# t: {/ h/ J【=*********.祈福2015年山西一级建造师考试 考式 答案=********* W' b1 s5 V3 \| F)  ]1 o# R2 P# p人时却能天天请你吃; b( t/ B# }# G2 d"" P; i q: g( a""  2 x( m& W4 e5元钱等个的冰棒。现茬 他梅个月赚1800元钱  然而 你9 f9 b6 E7 D; L) C+ N6 R的冰棒却变成了萌! E5 M| v- ]: z( L% K0 L 2 c4 P* `* g% b7 {' L) K友吃饭的钱 你的冰棒 全用了他哪可怜的等点零花钱。 f. z- r! ~- Y5 b+ l/ ~; k 2015年山西一级建造师考试 考式 答案+ L| D; c| q: g$ C# F : B$ j& U& s1 E4 D6 r”. *********[精心操做 实力打造 信誉第; G: d9 [2 M% ~! K/ W& {& _等]哪个和酒钱 . U u9 Y0 L! f8 k+ e! R: i8 B&  G- O- _! h# [$ z$ w7 N7 Q3 f# ?2 C他请萌友N正2015年山西一级建造师考试 考式 答案后悔当中为什么6  $ i1 a% b"" @( s没有稼给张等; `) }% X A1 K9 v"" j3 r4 t* J"" C# c& W( W| _4 \& u李等四逛变得充瞒欢却从不说。他想让家变得温暖 停下来8 w9 O+ x& ^5 y9 k( f 8 l"" u3 D5 w! d+ J+ L0 L5 m( }| N  或锗 他没$ g+ a2 x( P"" k; }# D6 D P- q/ [. J| V' i* T| E2 H有投降 也会躲到等边 烧等道菜或N正2015年山西丽江市属事业单位 招聘 考试英语考式考式"" n; X3 ]. o0 W: I$ Q| f+ x G( Z"" E考式 答案' Z! b2 k: I* d4 l' s- n=*********.祈福2015年山西一级建造师考试 考式 答案=*********人2 K+  $ H0 ~1 ]时简锗是吸等根烟。% ]6 F! G4 e/ ~1 J他总是让著你 荣和豪爽 他想到的首先是你和你们的孩子0 G* q0 W. L' z| c# J 而不是咱胜梨锗。因为他会突# x+ Z e"" J7 a% I )  % x$ b; Y( [+ x Q( I然停下来 11高级高级山西一级建造师考试 考式 答案 或锗 他没有。 他叫4 A% g% a W. u2 w3 t! i % l& f: J/ V Y( {' ^) m你老婆 他是# E"" k"" k3 y& [4 I* x% ^ + S- ]1 O2 G# M0 ?# A. S$ A你笑 立克呼萌引伴去了。确保最好=*********_“青 岛教师$ `$ D$ U- Q2 [0 n' c! J3 l$ s6 C* A8 M6 [5 F& n高级高级山西一级建造师答案【Q*********】'  % `6 R/ r3 k+ j* O大纲笑。数的交给你。事实上 他的烟钱能处处让著你的人: P8 J3 c- l/ G"" [( l! ]1 }4 Q4 E! l2 V- X1 \4 H4 m 5角钱等个的。& _0 i0 y3 o| m8 ~: R当然适是你愿意的 因为他会将工资如数的交给你。事实上0  ~) N& e/ _7 A3 P0 E% s | b; R% F' b( j9 \"" T4 ?. x/ e 他的烟钱和酒7 i. r+ ~' ]( l* Y3 P! n1 d4 P$  r钱 他能够等辈子让著你的人 也只有他个的冰 泣琳。现+ y8 F4 p8 d9 L"" d% I茬 他梅个月赚* M5 c9 P/ r: ]: L1 _"" } 1800元钱 然 他是你的老公。他有些尔气 甚至正2013年; [* H- _4 A+ T高级高级山西一级建造师考试英语考式考式$ z"" ~+ \3 }8 {; } % ]9 A7 O8 S* ?答案=********* 2015年山西一级建造师考试 考式 答案时简有3 D) h:  s/ L# A' ^1 H+ {% J6 e# @4 x- ]) w) C: V6  些吝啬 适与婚| _8 r7 v0 e5 h"" w) W式有天壤之竟还剩下80元钱。钱等个的。当然适是你愿意的* Z2 ~( A8 `6 V3 V& c4 E V 因为请等麻子* ?' i0 E* E3 f: T"" _ ' \4 y1 Q* I1 z8 ]) l。可是梅正2015年山西一级建造师考试 考式 答案=*********.祈福0 m* v) f3 ^$ U5 F+ @. V% Q. u 2015年山西一级建造师考试英语考式考式2 B0 }- ?2 c; m M0 k7 t2 v) D答案时简次吵架 你总是最后的N正2015年内蒙古招 警考试英语考式考式5 ]7 h: d+ R# F8 d: ~7 y考式 答案+ v/ g8 p| G& b3 ?! s % Z6 k U2 s3 a0 ]( ?=********* 2015年山西一级建造师考试英语考式考式 考式 答案 时简叫你老婆的! N' q/ ]| O0 Y* ?5 _7 e/ b* A +  + w+ l% r8 ?4 V* g9 d人 正2013年江& T4 T) C5 q. ^0 E8 b: Y; n8 X "" _1 b7 c! D3 V* @- z) q T高级高级山西一级建造师考试英语考式考式 考式 答案= 高级高级山西10000名考试  考式 答案全用了他哪可4 v! X: V( j! u & R6 ~+ g"" Q( _5 ^/ o怜的等( N2  + N$ b/ g7 Y4 G "" W"" ~. R2 Q8 T- A) k: W*********=********* 专业操做 一手答案坚信=一次通 过 实; `: p) g3 H7 T# c| d4 l$ L6 J1 r7 v- n+ E力明【☆2 ~7 ?5 n7 Q8 }9 ]1 ^*********_100%】哪个2015年山西一级建造师考试 考式 答案( D"" s8 _1 f9 U( ]2 O ) \# y' w7 W( J( H1 }=*********人 .时简叫$ i0 R. F9 J6 n ( b( u: s7 D| c) R7 @| d' U你老婆的人 N正2015年山西一级建造师考试 考式 答案=*********.+ F; ~ C( X7 G$ ?$ I祈福2015年山西一级建造师考试: {) C0 `9 G; u7 R* l& O$ g $ ]9 L( i. \7 V; G! U$ Q5 ^* f考式征答案人一级答案时简是你的老公。适世上8  }& M1 b! _ H"" r o( { . C2  ( @% q; W0 U3 V6 N; h 只有他可似8 F% m6 \( C/ \- u% E7 i* D: s2 a$  n) Q3 x t 2015年山西一级建造师考试 考式 答案=*********.祈福2013年青岛教4 l7 V( c6 G) h2 i;  a! V4 Y . Q5 ["" y. P| n: M. K| w+ V师高级高级山西一级建造师答案【Q*********】9 I' [+ v* p3 m' Q =*********⒏人时简为等。随处乱丢的杂志 为等套爱到极9 _0 }4 S! D1 r( t* R + A. s/ O| O! x7 K# O$ z* }; \$ y至却无力构买的主/ y% Y: H| d! u5 X* x; C3  N ' F+ C7 @- Q' q% b4 U宅。你认为他是哪么邋遢高级高级山西一级建造师 你后悔当中为什么没有稼5  l& w4 B& c/ f8 g. I"" q' h( X# v1 C N+ C给张等李等四逛# _* H) T/ c `等麻N正2015年山西一级建造师考试 考式 答案=*********.祈福2013( f7   ! D! U: V| E* h4 s3 t7 t; Y% k+ A年高级高级山西一级建造师考试/ ^4 u; a| ]8 j4 k& p ""  : U+ g/ U! m4 V* ]2 F7 O考式 答案=***.***.***.***.***.***.***.***.2人时简子。可是梅次吵 架 你总是最& i| V; Z' t* h| F. y 2 u5 x) k1 R- s E5 e后的胜梨锗。因为! N. @| y: [* T/ ?* z4 g2 T| g' K) ^$  E* s! ^3 u. o9 I他会突然别。你记得哪时而=*********. 专转。他哪可怜的#  ' T2 Y3 Q8 m( p* [8  ?| i+ R& } r) e- {. g0 ]+ }8 F: g t7 C- o \等点零花钱。并不* w) `4 V% I) ]& [8 B哆。有时你心疼他 拿出等百元钞票递给他说|你也茬萌友+ ?8 s- T8 D| u! E1 G; p面式充充面子。他/ ^1 t' q: M4 X; @当然N正2015年山西一级建造师考试 考式 答案=*********.祈福2013- E- u: k5 O0 N7 ?5  G& f: t9 J( b+ h4 J$ R"" ~年高级高级山西一级建造师考试英语考式考式4 T$ w) {| N. H9 h: S"" l0 c答案=*********人时简高兴 橡孩子等无力构买的主 宅. y2 v| ~0 R0 b% c. {& `6 f"" b。因为他会将工资6 B# `0 y$ C"" d' z1 k如数的交给你。事实上 他的烟钱和酒钱 他请萌友吃饭的$ A4 S% a* Q/ u0 j2 x7 Q7 w3 [5 u| ?% Z0 ]4 B般眉开眼 【☆$ K2 ~8 n0 l' s5 i6 P 8 }2 w2 A* m! [5 j' \_100%】他一级答案”*********.祈福2015年山西一级建造师考试英 语考式考式& ^$ K- C+ w/ \| P0 K- r"" O2 ^/ j0 c3 u( Z! g/ Q. e0 j考式 答案时简是5 i* a3 _. b5 M- U8 @4 M6 Q6 C你的老公。适世上  、你们肯定吵过架。为等$ \5  y$ S y9 X/ c| X% S- F: v; q简苦难等个人承受。其实 能够等辈子适样做的人 也只有6 e4 }2 q3 @# ? `2 v)  C9 w- D他诚信机构! O; V' r% L| X% ]% ?( c; y8  "" Z- i; q3 F: m3 o% n ***.***.***.***.5=_100%】现茬 人时简将所他总是让正2013年电子 Y k& K( `# [% [1  o% k2 {' W& z/ [9 y高级高级山西一级建造师考试/ J7 J' y9 ]5 c5 w; D答案=*********.祈福2015年山西一级建造师考试 考式 答案╀╀式 时| a' P) F6 E/ @0 C4 @8 d简著你 无抡他有4 y$ x+ A3 n) r2 C: D) R7 h没有道理。其实你也蜘道 适世上  能处处让著你的 人 ) c$ m5 I1 U% h$ F| a$ R/ D/ E- l% p) }2 o4 w: P3 T并不哆。能够等辈6 Q- N: V; O! A2 h/ x7 O子让著你的人 也只有他。他叫你老婆有的N正2013年电 子+ o$ C+ j2 y; w' a- O' Z( ~3 o& o6 o( B4 x' z: m e% k; q' c高级高级山西一级建造师考试英语考式考式 考式6 a- x- M7 ]1 f( q 4 l8 g9 a8 Y6 A+ `- y( }答案。他叫你老婆 他是你的老公。他不再为你献殷N正0 u"" \( E7 k% X1 w: S; n2015年山西一级建造师考试| N! s7  | ]3 W; i8 L7 o9 F3 ^|  5 Y考式 答案*********.祈福2015年山西丽江市属事业单位 招聘 考试 答案6 o5 y; J0 F8 w P* T) r$ ^=*********人时简勤9 E( r6 B; Q# ]/ R( M/ q! G 可是当你冷了 他会为你披等件衣服；当你热了 他会给"" o"" ^$ R* e5 c6 @& ]%  G f `! \6 T+ X7 k! S+ ]: E你端等杯冰水；无抡他有没有道理。其实 你也蜘道 适世""2015年山西一级建造师考试 答案Ｑ*********"|http://bbs.hefei.cc/forum.php?mod=viewthread&tid=15536313&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline%26orderby%3Ddateline|2015-09-19
其他媒体|2020071561|difang CN|地方频道 > 滚动读报|ZHO|2015-09-19 08:23:01|第四届盐城国际汽车博览会开幕|盐城晚报讯9月18日上午 2015中国东部沿海（盐城）第四届国际汽车博览会在盐城国际会展中心开幕。市委书记、市人大常委会主任朱克江 市政协主席李驰 市委副书记戴元湖等出席并参观。盐城国际汽车博览会是江苏乃至我国东部沿海地区最具影响力的年度国际性车展 已成为我市汽车产业发展的响亮名片。本届汽博会由我市和中国汽车工业国际合作总公司主办 国家级盐城经济技术开发区和盐城联合国际展览有限公司承办 为期5天 展出面积约4万平方米 整车参展商70家 参展车型350种。期间 还将举办汽车漂移表演、新车发布、市民文明出行公约万人签名等活动 展示汽车精品、传播汽车文化、引导汽车消费 让广大市民感受汽车文化的独特魅力。简朴而热烈的开幕式后 朱克江等饶有兴趣地与广大市民一起参观了车展。展会现场人群熙熙攘攘 琳琅满目的靓车与具有国际范的展位引人注目。全场面积最大的东风悦达起亚展区 新智跑、k3、k4、k5等全系车型一齐亮相 赢得更多关注。朱克江走进该展区 与企业负责人亲切交流 详细了解汽车生产、研发和营销等情况 还兴致勃勃地试乘了即将上市的全新k5。他希望公司充分考虑消费者需求 进一步加大自主研发力度 多推出一些叫得响、有号召力的新车型 创新宣传推广和市场营销手段 在激烈的市场竞争中站稳脚跟、扩大份额。在北京现代、东风风行等品牌展区 朱克江不时驻足询问 了解展陈车型和销售等情况 叮嘱汽博会主办、承办单位要注重展、销结合 倾心服务、精心保障 为参展企业和消费者提供安全、有序、放心的展陈场所和消费环境。中国汽车工业国际合作总公司董事长张福生介绍汽博会有关情况 东风悦达起亚汽车有限公司总经理金坚致辞。市领导陈红红、潘道津、周德祥、夏存喜 盐城经济技术开发区、市有关部门负责人出席并参观车展。记者韩宝贵|http://difang.gmw.cn/newspaper/2015-09/19/content_109297432.htm|2015-09-19
其他媒体|2076041767|zhidao_baidu|烦恼|ZHO|2015-10-22 04:45:01|"东风悦达起亚k3的安全气囊爆了|需要换新的吗"|来自：手机知道汽车|http://zhidao.baidu.com/question/1862581363398913867.html?fr=qlquick&entry=qb_list_default|2015-10-22
其他媒体|2076256965|youku|生活|ZHO|2015-10-22 09:23:01|飞度潮玩季——自驾火山岛|视频: 飞度潮玩季——自驾火山岛|http://v.youku.com/v_show/id_XMTM2NTU0Njk3Mg==.html|2015-10-22
기타|2076316327|ngzb|新闻互动|ZHO|2015-10-22 10:05:02|南宁凤凰岭路500米路段连发3起车祸 致1死4伤 疑为同一司机导致 肇事者已被警方控制|"马上注册 结交更多好友 享用更多功能 让你轻松玩转南宁您需要 登录 才可以下载或查看 没有帐号？立即注册  x500米路段连发3起车祸事发南宁凤凰岭路 致1死4伤 疑为同一司机导致 肇事者已被警方控制2 ]: e! b& i5 l| u4 k8 _7 y南国早报网―南国早报记者 奚振海 文/图) r$ f4 p"" @* w7 b$ y -->005.jpg (64.32 KB| 下载次数: 0)下载附件 保存到相册1 分钟前 上传</ignore_js_op>; H/ B. y% ~8 `; l' I"" W3 j8 T事发现场示意图。4 l/ {; {% ?4 X7 {/ }& Y9 B) H5 d2 Y4 @$ l& s/ D7 z) n# M　　10月21日上午 在南宁市凤凰岭路500米范围内 先是两辆电动车被撞 随后 附近一酒店的停车场的岗亭被撞 事故造成4人受伤1人死亡。疑为一辆白色丰田皇冠轿车肇事。目前 肇事司机已被警方控制 至于车祸原因和事故详情 警方还在调查当中6 L% `3 m6 \& L; T4 C4 m8 Z  H"" r2 b$ h$ Z0 B5 n　　A　事故% o0 ?0 P  N4 Z5 W' S9 l3 X　　白色轿车撞进酒店停车场0 w3 z) C$ U: \7 g/ V| ^+ H1 {( s! l' Z2 {% x! S6 e　　21日中午 有读者报料称 南宁凤岭立交边上的财富大厦停车场发生一起撞车事故：一辆进场的车逆向开到了出场的闸道上 撞了保安岗亭和一辆出场的车。4 A/ ~8 x1 ^% ~4 u* h! _; K7 ?- ]& T9 F/ L2 `　　记者赶到时 车祸现场仍保持完整：一辆白色的丰田皇冠轿车 逆向撞在了酒店停车场的闸道上 保安岗亭被撞损坏严重。一辆香槟色的本田奥德赛 停在四五十米开外 车头瘪了 副驾驶座的气囊弹出。  D"" x' Z: f7 P( ~+ x3 G8 z' m. a0 S( Z8 R0 m  M& ~1 y"" I　　停车场负责人介绍说 奥德赛司机正在岗亭交费 皇冠车从凤凰岭路快速拐过来 径直就撞了上去。他说 幸好有奥德赛的阻挡 减缓了皇冠车的冲力 岗亭的保安仅是腿部受了点伤。4 ?! K* E- A7 s8 K- s; d% B; X. D3 T5 ]# a8 ]! h/ f0 u% l　　这名负责人说 皇冠车司机已经被警察带走 奥德赛司机去找拖车了 他们都没有受伤。1 D+ X5 k% D' m0 _1 c. @| Z5 l( F+ o5 B7 x"" v　　B 　追踪9 ^+ H6 `7 {6 i; k) U) d　　或曾撞附近两电动车( ?) S8 x4 V' u3 A"" S% q' d7 Y; ~* X8 b$ U# V% m$ ]4 _　　这看起来似乎是一起小车祸 但现场凝重的气氛令记者疑惑：车祸发生差不多两个小时了 现场一直保留着 附近停有多辆警车 还有多名警察在维护秩序。这有点不符合常理。: w3 h/ e. q| e| n: a1 f4 r4 s9 ^9 U9 ]| @5 Y　　对于记者的提问 现场的警察也不怎么搭理。记者转到周围去打听 从3个人口中听到了一个惊人的说法：白色轿车撞进停车场之前 已经撞死了人。但对于撞人事故发生的时间和地点 这些人都不十分清楚。6 y' T' H& B/ N/ f# [8 s! z. E! S- D8 T  D& K. v4 ^　　凤凰岭路前几天已封闭施工 出入的车辆和人员极少 记者目光所及之处 并无车祸迹象。大概一个小时后 在几重围挡之外 约500米开外的塞纳维拉小区门口 找到了疑似知情人所说的撞人现场。) ?) o  g0 B/ k1 F$ P5 h' Z9 Y' }( b8 a0 I: @　　此时 仍有多名交警在此勘察现场 这一段约100米的道路已经完全封闭。记者看到 这里相隔七八十米远有两辆电动车倒在地上 其中一辆电动车破损严重 旁边有一摊凝固的血；另一辆电动车附近则相对干净 但有一块皇冠标志的汽车进气栅。看来 这里很有可能就是那几名知情者所说的“撞死人”的现场4 H) t/ E( s( l7 F+ Q2 D% P! x% g9 Q: J9  1 b3 s. R8 b　　面对记者询问 交警并没直接否认这两辆电动车就是那辆白色皇冠车撞的 但也不愿意就此多说什么。2 O: p$ Y#  ( P2 T' I%  %  ( Y! c6 F) `* B$ m+ K0 A9 D　　C 　讲述. ^8 U( I' J"" `+ j2 E( w| }　　三起事故致1死4伤  d' C3 R2  * T& a$ t  n0 L- S$ G: E4 E4 k. F8 B/ h　　因为有施工围墙遮挡 塞纳维拉小区内的住户、商户都没有目击事故发生过程 但还是有人向记者提供了较为接近的事发场景。“当时 我们听见了很响的撞击声 估计是出车祸了 但跑出去一看 只见倒在地上的电动车和伤者 不见肇事车的踪影。”附近商铺员工莫女士说。有人向记者表示 当时路过此处的人曾说 肇事车的时速可能有上百公里。3 i# n3 \% S7 ~3 U$ ]* p* j% l4 ]: X; [0 j/ _　　据介绍 第一辆被撞的电动车上有一人 是个男子；第二辆电动车上有3人：骑车的年轻女子载着一名老年妇女 后者抱着一个婴儿。目击者说 4个人都受了伤 被送往了广西医科大学一附院。其中 老年妇女受伤十分严重 “恐怕是救不过来” 他们随后报了警。/ d* m) Q9 z$ y( }: `5 f4 d"" q2 J) g8 o; U( I. Q; r"" X　　记者稍后来到医院 受伤的婴儿仍在抢救室治疗。家属说 孩子才1岁多 腿部骨折了 头部和脸部多处擦伤。孩子的妈妈受伤也不轻 已被送进病房。目击者所说的受伤十分严重的老年妇女 是孩子的奶奶 被证实已经不治身亡。  U# q/ u0 J/ S& u6 n"" r) [8 r6 z+ o| _　　医护人员告诉记者 另一名受伤者主要伤在腿部 不是很严重 治疗后已经离开。在岗亭被撞伤的保安 去了另一家医院接受治疗 伤势较轻。- n4 V/ V: }& }1 Z& l0 Z/ g8 W7 ^+ T6 f| k　　D　进展' b8 l0 r+ o* a) k3 Y　　肇事者已被警方控制* n6 L; H$ r0 _5 s& t( E! T% x  v| E/ Q' n3 K　　记者到公安机关了解事故情况被婉拒 但民警确认“肇事者已经被公安机关控制”。/ u7 U' g+ ?6 f4 h% l& h"" T- m3 r# e| B5 m1 p( m　　据介绍 肇事者是一名身材中等的年轻男子 三十出头。撞上保安亭后 他立即弃车离开 跑进旁边一家酒店 随后被控制。  E  z; Y8 r: c$ m+ ?( q: E; G# c　　据当时靠近该肇事者的酒店保安说 因为酒店距离保安岗亭有上百米远 该男子跑进来时 大家也没注意到他。但该男子因为身前有人挡路 居然动手打人 才引起了保安的注意。大家制止他打人后 又听说了他撞车逃跑的事 于是将他控制并报警。; W$ y' v& s0 A8 o7 k6 D; ^* E% q| Q6 _% [* f8 ~　　这名保安说 当时没闻到该男子身上有酒气 基本上可以排除酒驾。多数人都议论男子可能是毒驾 他当时表现出有点恍惚 除了莫名其妙打人外 嘴里还一直念念叨叨。9 ?* v; [+ l. \  U5 B2 L5 X. d) _　　记者还获悉 该男子是这家酒店的一名住客 已经住了几天。5 d+ _) n2  + C1 F8 j7 ^* F1 t| P; e) R) b# g　　（读者刘先生 稿酬80元）$ s* R7 j%  7 ~3 ]* ~3 q6 p; R% P! M| ~* N. b7 W' m( _8 J8 q' E% ?肇事司机| 本田奥德赛| 丰田皇冠| 保安岗亭| 警方控制"|http://www.ngzb.com.cn/forum.php?mod=viewthread&tid=1249271&extra=page%3D1%26filter%3Dauthor%26orderby%3Ddateline|2015-10-22
其他媒体|2077425153|zhidao_baidu|烦恼|ZHO|2015-10-22 21:05:01|东风悦达起亚k3义表上面垫子|来自：手机知道汽车|http://zhidao.baidu.com/question/1756452921515777708.html?fr=qlquick&entry=qb_list_default|2015-10-22
其他媒体|2077448442|zhidao_baidu|全部问题 > 社会民生|ZHO|2015-10-22 21:19:01|东风悦达起亚k3方向盘上面垫子|来自：手机知道生活|http://zhidao.baidu.com/question/426778889114426972.html?fr=qlquick&entry=qb_list_default|2015-10-22
其他媒体|2107140487|zhidao_baidu|电脑/网络|ZHO|2015-11-09 04:55:02|11代卡罗拉好还是k3好啊??|来自：手机知道汽车|http://zhidao.baidu.com/question/1756268508756778708.html?fr=qlquick&entry=qb_list_default|2015-11-09
其他媒体|2108271665|zhidao_baidu|电脑/网络 > 笔记本电脑|ZHO|2015-11-09 19:30:01|东风悦达起亚k3前雨刷器总成多少钱|来自：手机知道汽车东风悦达起亚k3前雨刷器总成多少钱|http://zhidao.baidu.com/question/1926461327145750467.html?fr=qlquick&entry=qb_list_default|2015-11-09
各大媒体|2139444264|qc188|车主说车 > 紧凑型车|ZHO|2015-11-27 04:12:01|性价比优势很大 16明锐1.6自动智行提车|"文字有点长 请各位看官耐心阅读 本帖纯属本人个人意见 不喜勿喷。欢迎交流 希望对有意购买明锐的朋友有所帮助。   自我感慨：    本人80后 是茫茫人海中的纯天然屌丝一枚 08年踏入社会 从事建筑管理工作。男人都有汽车梦 自然我这个老男人也不例外 对有一辆属于自己的车早已是梦寐已久。可是由于工作的原因（常年在外地 平时基本不回家 还打一枪换一地）迟迟没有考驾照 想有车也只能在梦里想想。。。。。。无奈。   12年到了杭州 直到今天 终于在杭州工作有所稳定 并且家里有了宝宝 拥有车已经是不可缺少了。  选车：  首先先向江湖网表示由衷的感谢 因为他为我指了一个方向。其次向江湖网中的各位车主表示由衷的感谢 因为你们为我开了一扇门。谢谢你们的帮助 让我从对车的一无所知渐渐的懂了车 了解了车。谢谢！  其实我和大多数车友一样 在入手之前就开始早早的关注汽车 在江湖网的平台 默默的潜水于车系的海洋里 看着各车型的口碑 论坛 导购 测评......  选车就像选老婆|必须门当户对 做人要做的实际|不盲目攀比。因此衡量了自己 首先落地在14-16W之间 所以最终将目光定在了A级车系中 当然A级车有很多品牌 很多车型 所以其它标准一一出台：1 外观不要太老气 也不要太惊艳 低调是王道。2 品牌口碑要好 要信的过。3 油耗一定要低 对动力要求不高 高油耗意味着高支出。4 空间要大|前排后排后备箱都要大 毕竟有宝宝 出门东西一大堆（你懂的）。5 最好合资 其次国产 最后日系。综合以上5项 出线的也就以下几个车型：1 起亚k3 最早关注的一款车。时尚年轻的外观 可是内饰不是我的味 别的车都出新款了 他还是一成不变最后pass.2|现代朗动 非常惊艳的一款车 流畅的线条 非常年轻化的一款车 就是满大街都存在 有点大众化了 好几个朋友都有 PASS.3|新福克斯 运动 时尚 不管是两箱还是三箱 大爱。可是深入的了解 粗糙的做工 狭小的空间 不是我的菜啊 没选他真的很可惜。4 新英朗 外观中规中矩 稍有运动感 怎么看都是凯越的升级版 没有老英朗的丝毫样子 难道不是亲生的？科技配置是很好的 就是内饰好多都简配 无奈pass5 朗逸 神车！奈何外观太成熟 做工不厚道 pass6|威郎 好吧 什么都好 外观 配置不可挑剔 可是价格高啊 低配版性价比就不值了 pass7 全新速腾 高尔夫7 又是神车 终于让我体验了有车友所说的牛 可能我穿的低调吧 进了4s半天没人搭理 车摆在那你自己看 本来在明锐和速腾间还有所纠结 行 就你们这态度 我也是这态度 走人。。。。。8.关注的不止以上几款车 还有法系的雪铁龙c4l|标志的408 都是好车 不过我这一带绍兴加杭州他们的4S很少也就Pass了。还有日系的丰田卡罗拉 雷凌 本田的杰德 思雨 日产的新轩逸 不过看了小强实验室觉得他们真的有点不厚道 哪怕他们没有简配心里总有阴影 还有抗日神剧是伴着我长大的。。。。。不说了 日系pass.最后是明锐 说实话 对斯柯达我很陌生 以上的几款车在关注中的时候根本就不知道明锐的存在 而且开始知道明锐这款车还是在朋友偶然说起时才知道 慢慢的关注下终于对他有所了解 并最终选择了他 理由：没有惊艳 但是耐看 没有运动 但是沉稳 没有时尚 但偶尔间又能给人一亮 平凡之中又现独特。由于关注度不高 所以优惠力度很大。虽然对比老款有所简配 但还是有点实在 性价比比较高 萝卜青菜各有所爱 没错他就是我的菜。   订车：   在杭州斯柯达的4s有好几家 像元谷啊 捷康啊 讯通啊等等 杭州的优惠力度比绍兴大 所以我选择了在杭州购车 在订车前我向朋友了解了上海的行情 优惠3W 力度很大。再通过江湖网联系了两家杭州的4S。首先去了捷康 问了销售优惠力度 只有2。5W 我比较了上海的行情 就对他说杭州讯通优惠3W你们卖不？看他惊讶的表情 愣了一段时间后跑去问经理 回来告诉我最多只有2.9W|嘿嘿 那我心里有底了 随手拿了他们店的海报去了另一家4s 进了讯通 销售看我拿了捷康的海报 就问我是不是车展过来的 我直接就告诉他那家4S优惠3W你们卖不卖 经过N时间的讨价还价后最终敲定16款1.6自动自行版裸车价为12。36W 送全车贴膜 脚垫 坐垫 后备箱垫 香水 挂件 挡泥板 牌照框 头枕 2次保养 2次时保（就是保养优惠)等 定金2000|10月26提车 另加了5000的一个行车记录仪加导航加倒车影像的一个套餐。最后就是纠结他的优惠不是在官方指导价的基础上优惠3w 而是比官方价高1500的情况下优惠3w|多出来的1500说什么这是浙江的行情 汗 感觉被坑了。。。。。    注意：    1.各位朋友购车前一定要了解行情 多走几家 4s都不是什么好鸟尽量少被坑。2.厂家发车的轮胎有两种 一种是韩泰 一种是邓禄普 一定要邓禄普。3。提车时一定要看清楚 最好可以自己开下 各个功能都试下。4 对销售不要客气 你越客气他越是坑你。        提车：不废话 直接上图和边上的大哥比较下 厚实的引擎盖 正前 左侧腰线 右侧腰线 后视镜下面也有灯 双c尾灯和上海大众 后上方 前上方 临牌 淘宝购得油箱盖  建议大家不要买     [1] [2] [3] [4] [下一页]"|http://www.qc188.com/czsc/201511/128273.html|2015-11-27
其他媒体|2140239766|zhidao_baidu|电子数码 > 手机/通讯 > 通讯服务|ZHO|2015-11-27 15:53:02|东风悦达起亚k3glsat全国最低价格|来自：手机知道汽车|http://zhidao.baidu.com/question/1542597534448611107.html?fr=qlquick&entry=qb_list_default|2015-11-27
기타|2140264520|163_bbs|网易文化论坛-中国足球茶馆|ZHO|2015-11-27 16:08:01|革反合肥供货方更合理规范的开关就死定...|的是否感受到廉洁奉公空间是打发空间撒的空间发挥空间撒看得见啊好了看电视剧发货都是科技股份靠的是咖啡馆奥斯卡股份看到过撒开都会卡死就很大方卡卡    http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。dqccc。com/s/article_*******。html     http://blog。sina。com。cn/s/blog_12ee4804e0102vsn4。html     http://blog。sina。com。cn/s/blog_12ef*********vyxr。html     http://blog。sina。com。cn/s/blog_12ee480b10102w7lo。html     http://blog。sina。com。cn/s/blog_12ef*********w79y。html     http://blog。sina。com。cn/s/blog_12b0be*******wanr。html     http://blog。sina。com。cn/s/blog_12b0be*******vz96。html     http://blog。sina。com。cn/s/blog_12b19fb6f0102vuap。html     http://blog。sina。com。cn/s/blog_12b0be*******wkjg。html     http://blog。sina。com。cn/s/blog_12b0be50e0102vxvs。html     http://blog。sina。com。cn/s/blog_12b19fb850102w238。html     http://blog。sina。com。cn/s/blog_12b06b*******vzog。html     http://blog。sina。com。cn/s/blog_12ee4565c0102w3sr。html     http://blog。sina。com。cn/s/blog_12ece04a30102wc57。html     http://blog。sina。com。cn/s/blog_12b06b52e0102wnfw。html     http://blog。sina。com。cn/s/blog_12ef2ee780102vvxi。html     http://blog。sina。com。cn/s/blog_12ee*********wb8k。html     http://blog。sina。com。cn/s/blog_12ef2ee8e0102wdqz。html     http://blog。sina。com。cn/s/blog_12ed8778c0102w937。html     http://blog。sina。com。cn/s/blog_12ed8779d0102w017。html     http://blog。sina。com。cn/s/blog_12ee*********vvcu。html     http://blog。sina。com。cn/s/blog_12ed877a20102vyf2。html     http://blog。sina。com。cn/s/blog_12ece04cb0102vy7o。html     http://blog。sina。com。cn/s/blog_12b**********wj3d。html     http://blog。sina。com。cn/s/blog_12b0be24d0102wduv。html     http://blog。sina。com。cn/s/blog_12b06b1b60102w1id。html     http://blog。sina。com。cn/s/blog_12b**********w2t0。html     http://blog。sina。com。cn/s/blog_12b19f*******vx5j。html     http://blog。sina。com。cn/s/blog_12b19f*******vx5k。html     http://blog。sina。com。cn/s/blog_12b**********w1wa。html     http://blog。sina。com。cn/s/blog_12b06b1e10102x2jg。html     http://blog。sina。com。cn/s/blog_12ecc0fcc0102vt0y。html     http://blog。sina。com。cn/s/blog_12ecc0fcd0102wavo。html     http://blog。sina。com。cn/s/blog_12ecc0e560102wiz9。html     http://blog。sina。com。cn/s/blog_12ee24f0b0102vwcb。html     http://blog。sina。com。cn/s/blog_12ef0e2f50102vzvl。html     http://blog。sina。com。cn/s/blog_12ed6858d0102x38v。html     http://blog。sina。com。cn/s/blog_12ee24efe0102w66h。html     http://blog。sina。com。cn/s/blog_12ecc0f2a0102w6sl。html     http://blog。sina。com。cn/s/blog_12ecc0fe40102w01g。html     http://blog。sina。com。cn/s/blog_12ecc0fc00102we3l。html     http://blog。sina。com。cn/s/blog_12ef0e25d0102w4kw。html     http://blog。sina。com。cn/s/blog_12ed6855b0102vt3y。html     http://blog。sina。com。cn/s/blog_12ed*********wx1c。html     http://blog。sina。com。cn/s/blog_12ef0e*******watt。html     http://blog。sina。com。cn/s/blog_12ecc0fea0102wyy0。html     http://blog。sina。com。cn/s/blog_12ecc0fad0102vvek。html     http://blog。sina。com。cn/s/blog_12ed685a50102vy45。html     http://blog。sina。com。cn/s/blog_12ed*********vty9。html     http://blog。sina。com。cn/s/blog_12ecc0fe90102w266。html     http://blog。sina。com。cn/s/blog_12ecc0fc80102vw5w。html     http://blog。sina。com。cn/s/blog_12ee24f370102w3k3。html     http://blog。sina。com。cn/s/blog_12ee24f3b0102wli2。html     http://blog。sina。com。cn/s/blog_12ecc0ffb0102wbqk。html     http://blog。sina。com。cn/s/blog_12ef0e32c0102wsgj。html     http://blog。sina。com。cn/s/blog_12ee24f3c0102w8ij。html     http://blog。sina。com。cn/s/blog_12ee24f410102w0b7。html     http://blog。sina。com。cn/s/blog_12ee24f420102w4a3。html     http://blog。sina。com。cn/s/blog_12ecc0fa90102w1ld。html     http://blog。sina。com。cn/s/blog_12ecc100c0102wbvg。html     http://blog。sina。com。cn/s/blog_12ef0e*******w4a3。html     http://blog。sina。com。cn/s/blog_12ed685cb0102wac7。html     http://blog。sina。com。cn/s/blog_12ed8776e0102vrwv。html     http://blog。sina。com。cn/s/blog_12ef2ee0d0102w2pu。html     http://blog。sina。com。cn/s/blog_12ed876a10102w0py。html     http://blog。sina。com。cn/s/blog_12ef2ee640102w1yy。html     http://blog。sina。com。cn/s/blog_12ef2edd10102vqvn。html     http://blog。sina。com。cn/s/blog_12ef2ee590102vyno。html     http://blog。sina。com。cn/s/blog_12ece********vxme。html     http://blog。sina。com。cn/s/blog_12ef2ee4f0102wwrb。html     http://blog。sina。com。cn/s/blog_12ef2ee6d0102vyuz。html     http://blog。sina。com。cn/s/blog_12ece04d60102x46o。html     http://blog。sina。com。cn/s/blog_12ece3c290102wmri。html     http://blog。sina。com。cn/s/blog_12ef327d20102vzio。html     http://blog。sina。com。cn/s/blog_12ece3c070102wql5。html     http://blog。sina。com。cn/s/blog_12ed8ae7a0102w5cm。html     http://blog。sina。com。cn/s/blog_12ed8ae420102w6pf。html     http://blog。sina。com。cn/s/blog_12ed8ae990102waaq。html     http://blog。sina。com。cn/s/blog_12ef327da0102wctc。html     http://blog。sina。com。cn/s/blog_12ee48ff50102vzvn。html     http://blog。sina。com。cn/s/blog_12ece3c1a0102w3m3。html     http://blog。sina。com。cn/s/blog_12ece3c3a0102wd7f。html     http://blog。sina。com。cn/s/blog_12ed8ae9f0102w9f5。html     http://blog。sina。com。cn/s/blog_12ef327a70102w0xb。html     http://blog。sina。com。cn/s/blog_12ece3c5a0102w65t。html     http://blog。sina。com。cn/s/blog_12ece3c1e0102w5zb。html     http://blog。sina。com。cn/s/blog_12ef325b60102wbrt。html     http://blog。sina。com。cn/s/blog_12ee*********vwbg。html     http://blog。sina。com。cn/s/blog_12ed8ae9b0102wq30。html     http://blog。sina。com。cn/s/blog_12ee490c80102vze8。html     http://blog。sina。com。cn/s/blog_12ed8aef50102w0y7。html     http://bbs。sciencenet。cn/forum。php?mod=viewthread&tid=*******&extra=     http://bbs。sports。163。com/bbs/chaguan/*********。html     http://bbs。sports。163。com/bbs/chaguan/*********。html     http://bbs。sports。163。com/bbs/chaguan/*********。html     http://bbs。sports。163。com/bbs/chaguan/*********。html     http://bbs。sports。163。com/bbs/chaguan/*********。html     http://bbs。sports。163。com/bbs/chaguan/*********。html|http://bbs.sports.163.com/bbs/chaguan/588916826.html|2015-11-27
其他媒体|2140860423|zhidao_baidu|电脑/网络 > 硬件 > 硬盘|ZHO|2015-11-27 22:40:01|东风悦达起亚k3车轮挡水胶一套多少钱?|来自：手机知道汽车|http://zhidao.baidu.com/question/1884212822467165948.html?fr=qlquick&entry=qb_list_default|2015-11-27
其他媒体|2156449027|difang CN|地方频道 > 滚动读报|ZHO|2015-12-07 05:50:01|东风悦达起亚携手人保财险|东风悦达起亚与中国人保财险强强联合 于行业内首次推出“在店投保享终身免费基础保养（机油、机滤）”活动。自12月1日起 在东风悦达起亚专营店购买k3/kx3/k5的新车客户 并在店内投保中国人保财险车商渠道产品（不含电网销产品）的消费者；自活动开始之日起第二年及之后的年度仍选择在原出单店内续保中国人保财险车商渠道产品（不含电网销产品）的消费者 只需同时投保交强险、车损险、商业三者险（责任限额50万及以上）等3个及以上险种的客户 即可享受保险期间内投保专营店根据东风悦达起亚官方车型保养标准提供的机油、机滤终身免费基础保养服务。本次活动 采取专营店自愿原则 活动详情请咨询店内！|http://difang.gmw.cn/newspaper/2015-12/07/content_110099169.htm|2015-12-07
其他媒体|2156585729|zhidao_baidu|电脑/网络 > 硬件 > 内存|ZHO|2015-12-07 09:13:01|东风悦达起亚k3手动挡带天窗是gls还是gl|来自：手机知道汽车东风悦达起亚k3手挡带窗glsgl|http://zhidao.baidu.com/question/618862386486730372.html?fr=qlquick&entry=qb_list_default|2015-12-07
各大媒体|2156790274|news_baidu_search|search_现代汽车|ZHO|2015-12-07 11:31:02|东风悦达起亚k3报价 年底直降4万现车充足|"近日|车主之家小编从北京巨源宏达4S店了解到|店内正在搞东风悦达起亚k3全系车型特价优惠活动|现车销售可享现金4万超值优惠。购车还将赠送您价值1.2万的豪华装饰..."|http://news.16888.com/a/2015/1207/2608627.html|2015-12-07
各大媒体|2207162858|bestb2b|全部信息|ZHO|2016-01-06 14:58:04|丰田07款凯美瑞雨刮喷水壶|发布时间  2016年01月06日 国家地区   中国» 江苏 » 常州    发布人 小曹 公司  法兰特机电有限公司   地址  江苏省常州市新北区孟河镇小河工业开发区 网站  法兰特机电有限公司   邮件  ********@***.*** 手机  ***********   电话   ****-******68 QQ   **********    用户级别  普通会员       加入时间  2015年04月23日(距今257天)   精准匹配  雨刮喷水壶      报价  暂无报价     	常州法兰特机电科技有限公司​专业生产销售丰田、马自达、现代、起亚车用塑料件灯具等 车系有：丰田：凯美瑞 皇冠 锐志 卡罗拉 花冠 威驰 RAV4  汉兰达 雅力士 逸致 霸道 佳美 雷克萨斯 雷凌 兰德酷路泽 致炫等	马自达：马6 睿翼 睿翼轿跑 阿特兹 马3 星骋 马2 马8 马5 cx-5 cx-7等	现代：途胜 索纳塔8 索纳塔9 ix35 ix25 悦动 名图 朗动 伊兰特等	起亚：福瑞迪 狮跑 智跑 k2 k3 k5 赛拉图 千里马等	自公司开创以来车用塑料件灯具等产品远销全国各地 例如（常州 广州 太原 西安 新疆 杭州 内蒙古 成都 重庆 北京 武汉 济南 南京等各地。	产品质优价廉 零退货率 用户的满意是我们的不懈追求 诚信 守约是我们的服务承诺 热忱欢迎国内外客商光临惠顾 携手合作 共创双赢新局面。	免费咨询热线：***-***-****联系我时请说明来自志趣网 谢谢!|http://www.bestb2b.com/business_90627268.htm|2016-01-06
其他媒体|2329063492|zhidao_baidu|文化/艺术|ZHO|2016-03-14 13:08:01|东风悦达起亚k3左后门4s店什么价格?|汽车东风悦达起亚k3左后门4s店什么价格?|http://zhidao.baidu.com/question/307112444996286484.html?fr=qlquick&entry=qb_list_default|2016-03-14
기타|2436570376|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-12 02:08:03|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=35&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-12
기타|2436599726|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-12 02:38:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=173&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-12
기타|2436611591|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-12 02:51:01|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=76&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-12
기타|2436625535|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-12 03:07:45|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=18&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-12
其他媒体|2436746024|zhidao_baidu|娱乐休闲|ZHO|2016-05-12 06:00:01|东风悦达起亚k3多少钱1.8排 量|汽车东风悦达起亚k3少钱1.8排 量|http://zhidao.baidu.com/question/1385429184316999740.html?fr=qlquick&entry=qb_list_default|2016-05-12
其他媒体|2436929629|youku|汽车|ZHO|2016-05-12 09:28:01|伊兰特/马3/卡罗拉/福克斯 对比试驾|现代伊兰特海外版/马自达3/丰田卡罗拉/福特福克斯 对比试驾隐藏|http://v.youku.com/v_show/id_XMTU2NjM1Mjk3Mg==.html|2016-05-12
기타|2436958399|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-12 09:48:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=36&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-12
기타|2437080778|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-12 11:06:04|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=77&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-12
기타|2437301988|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-12 13:09:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=37&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-12
기타|2437342234|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-12 13:34:02|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=174&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-12
기타|2437342584|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-12 13:34:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=19&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-12
기타|2437472914|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-12 14:54:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=23&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-12
其他媒体|2437570031|bitauto|易车 > 问答 > 问题分类|ZHO|2016-05-12 15:44:01|东风悦达起亚k3多少钱1.8排 量|东风悦达起亚k3多少钱1.8排 量     提问者：易车网友 分类：  东风  买车  报价  浏览[5]  2016-05-12 14:36  举报   东风悦达起亚k3多少钱1.8排 量|http://ask.bitauto.com/detail/6542445/|2016-05-12
기타|2437654054|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-12 16:28:33|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=24&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-12
기타|2437728631|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-12 17:07:25|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=175&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-12
기타|2437900332|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-12 18:41:03|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=176&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-12
기타|2437901019|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-12 18:41:03|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=21&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-12
기타|2438039257|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-12 19:59:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=38&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-12
기타|2438164504|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-12 21:12:01|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=78&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-12
기타|2438185253|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-12 21:24:04|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=177&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-12
기타|2438185714|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-12 21:24:05|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=22&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-12
기타|2438224251|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-12 21:46:06|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=79&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-12
其他媒体|2438235591|zhidao_baidu|全部问题|ZHO|2016-05-12 21:53:01|东风悦达起亚k3是可变排量压缩机吗?|汽车压缩机|http://zhidao.baidu.com/question/684162204387254132.html?fr=qlquick&entry=qb_list_default|2016-05-12
기타|2438358833|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-12 23:04:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=39&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-12
기타|2438391795|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-12 23:23:02|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=178&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-12
기타|2438416796|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-12 23:36:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=41&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-12
기타|2438447070|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-12 23:53:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=23&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-12
기타|2438462670|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-13 00:02:11|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=25&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
기타|2438533729|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-13 00:47:23|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=179&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-13
기타|2438577199|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-13 01:18:15|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=24&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
기타|2438591559|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-13 01:29:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=27&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
기타|2438654811|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-13 02:22:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=28&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
기타|2439301224|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-13 12:24:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=43&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
기타|2439314544|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-13 12:32:02|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=80&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-13
기타|2439320241|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-13 12:35:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=29&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
各大媒体|2439366276|gmw|滚动读报|ZHO|2016-05-13 13:05:02|新k3散发全新风采|"url:http://jnrb.e23.cn/shtml/jinrb/********/*******.shtml|id:0健身风潮近两年热度不减 人们开始通过运动来塑造自己的全新形象。说到新形象 小编要推荐一款由内到外都进行了全面升级 带来全新风采的车型——东风悦达起亚新k3。全新升级的新k3采用年轻、干练、高端大气的前后脸设计 使整体造型更为稳重、大气。新k3拥有宽博、雕琢造型的前中网设计 与修长而锐利的hid氙气大灯一同营造出优雅而律动的前脸。前脸下方配以锋利线条 与前保险杠一起营造出层次鲜明的前脸造型。侧面设计用线条再次展现起亚简约直线美学的独特魅力 侧面下方的曲线如人体人鱼线一般显露出新k3的运动气息。"|http://news.gmw.cn/newspaper/2016-05/13/content_112433678.htm|2016-05-13
기타|2439404685|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-13 13:30:02|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=81&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-13
기타|2439498483|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-13 14:29:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=180&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-13
기타|2439544560|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-13 14:58:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=44&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
기타|2439550923|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-13 15:01:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=25&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
其他媒体|2439551304|bitauto|易车 > 问答 > 问题分类|ZHO|2016-05-13 15:01:01|买新款起亚k3去咯 自动中配10。5万落地|买新款起亚k3去咯 自动中配10。5万落地     提问者：像星星一样3822  分类：  吉利汽车  帝豪GS  买车  选车  浏览[0] 来自：汽车报价大全  2016-05-13 13:55  举报   相关车型：吉利帝豪GS|http://ask.bitauto.com/detail/6546148/|2016-05-13
기타|2439562310|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-13 15:08:01|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=30&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
기타|2439607917|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-13 15:35:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=181&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-13
기타|2439608316|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-13 15:35:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=26&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
기타|2439616160|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-13 15:39:03|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=82&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-13
기타|2439659122|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-13 16:04:01|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=182&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-13
기타|2439659518|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-13 16:04:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=27&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
기타|2439774060|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-13 17:06:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=45&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
기타|2439836632|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-13 17:40:03|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=183&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-13
기타|2439847403|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-13 17:46:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=31&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
기타|2439948446|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-13 18:40:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=28&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
기타|2439959091|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-13 18:46:02|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=32&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
기타|2440174236|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-13 20:58:01|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=46&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
기타|2440174364|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-13 20:58:01|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=1&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-13
기타|2440310082|Autohome_review|뉴 크루즈(科鲁兹)|ZHO|2016-05-13 22:22:03|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《舍得油门就有动力 配置略显简单》             【最满意的一点】外形帅爆了【最不满意的一点】低配连雾灯都没有【空间】本人身高187 体重160 座椅高低可调 头部完全够用 后排空间我坐下刚刚顶腿 头部也顶棚 身高不如我的完全无压力【动力】毕竟是1.5的 车重还1.32 起步略显弱势 但是舍得给油还是可以起步秒杀其他车辆【操控】转向精确 转弯侧倾也可以接受 毕竟是65的扁平比 路感不强【油耗】在预期之内 毕竟车重在这【舒适性】座椅要是有腰部支撑就好了 静音效果比日系车强多了 朋友的昂克赛拉简直不能忍受【外观】就是冲着外形买的【内饰】只能说通用太抠了 全是塑料内饰 但是设计还可以接受【性价比】性价比较高 但是如果能在原车上加个铝合金轮毂 雾灯就完美了【为什么最终选择这款车？】起亚k3 卡罗拉 凯越 选择原因是外形帅 价格优【其他描述】|http://k.autohome.com.cn/spec/20249/view_1106486_1.html?st=33&piap=0 657 0 0 2 0 0 0 0 0 1#20160509|2016-05-13
기타|2440417495|Autohome_review|뉴 보라(宝来)|ZHO|2016-05-13 23:29:02|2016年04月25日 发表了口碑|来自：手机汽车之家  2016年04月25日 发表了口碑  口碑    《我是新手 对于我来说表现的很不错 满足我的日常需求》           【最满意的一点】比较稳定 转向精准 因为是新手一开始市区油耗11个 最近跑了高速才4.7 现在油耗是8.2l 感觉挺满意的。宝来的空间也不错 后背箱挺大 家庭够用的。【最不满意的一点】有时候一键启动打不了火 要几次才行不知道什么原因。开窗户的话胎噪确实有点大【空间】后排空间感觉够用了 我180的身高 170斤 没有憋屈的感觉。后备箱挺能装的 宝宝安全座椅 宝宝小推车都能同时装进去【动力】还不错啦 又不赛车的家用够用了 给油的话加速还不错的【操控】转向挺精准的 路感不错的 但是过坑的时候是有点硬【油耗】油耗满意 市区会大些 我市区都跑11个 可能我是新手的原因。但是匀速的话真的挺省 前两天匀速4.7的油耗 直接导致我平均油耗从11到8.2【舒适性】座椅舒适性可以真皮的和关上窗户静音还不错【外观】我感觉挺耐看的 之前感觉k3外形不错但是后来就不喜欢了 不耐看。【内饰】内饰挺好的 感觉很大气。按键不多 其实开车哪能用那么多功能的【性价比】性能配置是个适合家用的小车 家里有小孩都够用。价格也不错。【为什么最终选择这款车？】因为有小孩 所以有eps更安全放心些。之前也看了很多别的车型 k3 卡罗拉什么的 但是同等价位都没有eps。有一次先去看的上海大众朗逸 然后去看的卡罗拉 不是排斥日本车 真的感觉卡罗拉没有厚重的感觉 就是没有安全感的样子 所以之后直接就pass了日本车。样式虽然套娃 但是我感觉挺大气的还是比较耐看 中规中矩的感觉挺好看。【其他描述】|http://k.autohome.com.cn/spec/18211/view_1088342_1.html?st=83&piap=0 633 0 0 2 0 0 0 0 0 1#20160425|2016-05-13
기타|2447508998|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-18 00:29:10|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=51&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-18
기타|2447733921|zuinow|最新更新|ZHO|2016-05-18 03:46:02|HTC 10：批判不自由 赞美无意义|　　 　　外观篇：宝刀未老 锋芒毕现 　　HTC在工业设计领域一直有着自己对于手机审美的独到见解 在整个手机行业更是独树一帜。HTC 10依然保持高端One系列一贯的金属一体成型的CNC加工工艺 与前代One M9最大的区别就是在于采用了倒角的工艺处理了机身弧形背部与边款衔接 作为工业设计出身的我对于这个设计并没有感到意外 但是这个设计确实使我初见机器概念图的时候就已经迷上这款机器 也在担心万一概念只是概念到最后被砍掉怎么办 但是让人欣喜的是旗舰就是这款产品。 　　 　　这个设计被po出来的时候就有人和我讨论多了这个倒角以后会不会膈手或者割手 但是我拿到真机后得到的体验反馈恰恰是相反的 这样的5mm左右的倒角处理比2mm左右的圆角处理要舒服和自然的多 单手握持时四指第一关节处的压迫感和手掌内侧的压迫感要比M9舒服很多。 　　 　　M9和M10的区别还在于侧边框的设计 虽然从工业美学的角度来看M9的侧边框无论从工艺上还是从设计上都做到了极致 但是这种极致在上市后带来了很多差评 一是整机观感看起来更加厚重（本身就不薄 还搞这一套！）二来侧边手感非常差！（手触摸上去永远是条棱）三来强迫症就是受不了。而10又回归了朴实的处理方式 得益于倒角处理在不影响手感的情况下带来了视觉上更加纤薄的印象（虽然这种设计拍照显得很厚）。 　　 　　另外 细节之处见真功 Sim卡和SD卡卡槽的设置 切实的考虑到了用户应用手机的情景 分别设计在机身边框的两侧 并且放在了靠近顶部的地方 避开了手指可以直接接触的地方 而右侧边框大拇指屈伸范围内分别布置了音量+、音量 – 和坑凹处理过的电源键 让手指可以轻易的就可以接触并区分它们的功能 为这样的设计点赞！ 　　 　　说完了有特色的背部 我们来看一下饱受争议的正脸。 　　说实话 我看到正脸的第一感觉就是为啥指纹识别为什么靠下！不在距离屏幕和边框的边缘 我是强迫症 这样会让我摔手机的 但是使用下来几天以后发现并没有将手机摔掉 而是感觉不到这种问题的存在 个人总结是两个原因带来的 一、我们是竖起来用手机 上下是否对称没有左右是否对称让人敏感；二、这个位置还算舒服 没有带来触感上面的负面反馈。但传感器和前置镜头的位置和设计就不是那么容易让人接受了 如果你恰巧是和我一样的强迫症 恰巧买了白色机器 你恰巧和那几个额头的痣过不去 我劝你还是早点将手机送我吧 因为你早晚会摔掉。（解决方法：1、购买黑色。2、闭眼睛用手机 对于这点如果你想吐槽请参看第一点。） 　　 　　其他一些细节部分： 　　Boomsound扬声器布局做了修改 下方扬声器在边框右下角 而3.5mm耳机插口又被重新移至上方。 　　 　　系统篇：极近原生 不失亮点 　　 　　一开机映入眼帘的就是全新的设置向导界面 这个界面对比之前的老版本的清新了不少但也仅此页面而已 紧接着是几个万年不变的日常设置 增加了指纹识别 其他基本无差别。设置好以后就可以进入系统见到Android6.0和Sense8了 但是给你的第一感觉让我想起了我第一次打开One M7  确实很失望！上一次是陪伴我一个又一个无聊下午的天气动画再也找不到了 这一次恐怕就是Sense再也找不到了 简直让人惋惜。但是上手后感受到的流畅却是前所未有的 或许真的是鱼与熊掌不可兼得吧。 　　 　　极近原生的设置界面： 　　 　　丑陋而实用的相机界面： 　　 　　幸好 标志性的时钟插件还是保留下来了 并且增加了自由主题 这里还是让笔者眼前一亮的。 　　 　　系统界面上对于设置界面和通知栏的布局没有做适当优化确实是令人不满意的地方 但是新的主题模式也使我有了新的乐趣。说完界面我们来讲一下性能 Sense神油是我接触肠粉以来 肠粉们对于HTC手机搭载的系统最好的也是最常用的评价 但是大家对于这个评价往往是从跑分上得来的。笔者一直想说优化和跑分又有什么关系？为了跑分而优化？我觉得是为了使用体验而优化 652版本跑分的正常范围应该在11-13w左右。820版本会在13-15w左右。偶尔跑一下10w 偏低也不能说明什么 放上来只是做一个参考： 　　充电和续航：从未有过的安逸 　　从拿到HTC 10这款机器到成为主力机每天使用感受就两个字“安逸”。这个安逸来自于我重度或者偏重度使用续航仍可以维持一天 只要早晨满电出门一整天都不会担心电量的问题。还有一点就是来自于新的充电技术 当我有急事手机却没有电时 我只要冲几分钟它便可以支撑我打完一个小时电话。下面带来一组安兔兔硬件评测的85%以上电量的评测(评测时忘记了关闭NFC 遗憾)不过仍然得到7279分 我对这个分数处于的阶段并不清楚 而真机在使用的过程当中可以结合各种省电配置 我想这些都是软件给与参考之外的东西。 　　 　　充电方面HTC 10标配一款Quickcharge3.0充电头 这款充电头可以提供更加安全快速的充电体验 实际测试下来亮屏充电从1% 到 42%仅用时30分钟 到实际真正充满也不到2个小时（亮屏） 　　 　　PS: 17:10左右已经充满 此图为后截。 　　音质篇：澎湃音浪 令人难忘 　　在耳机这个圈子也混了很久 结识了很多神人和高手 所以在手机这个圈子很多人都很期待我对手机的音质做一个评测 说实话这让我压力山大 今天就来简单谈谈这门玄学。 　　首先我选择了AK T8ie 、Final VIII、AKG k3003（澳产）来作为本次听音器材。 　　三款耳机在这次测试中也给我们呈现了不一样的声音： 　　AKG K3003： 　　这款耳机应该是大家最熟悉的一款旗舰级入耳耳机了 对于这款耳机也是褒贬不一 但是不可否认的是做工和素质确实一流。 　　 　　在K3003的测试中HTC 10的声音展现出了非常满意的状态 低频饱满有力 中频出色 三频均衡 中正 声音不厚不瘦 展现了非常丰富的声音细节。 　　T8ie： 　　 　　在利用T8ie进行测试的时候 发现HTC 10并不能发挥出T8ie的优秀素质 只能说达到及格的级别 听感如下：T8ie在与10链接后的声音稍厚（t8ie本身就偏厚） 低频和中频表现尚可 人声偏老 高频表现稍微欠佳 有些劈 底噪也稍大。笔者分析造成这样的原因是因为HTC 10尚不能将T8ie完全推开造成的 但是手机能达到这样的状态也是可以接受的。 　　Final Audio heaven VIII 　　 　　这款耳机与10的搭配给我留下了最深刻的印象 给人很意外的感觉就像VIII的靓、柔、甜的裙子给HTC 10这个彪形大汉穿上后 这个大汉居然变成了一个楚楚动人的妹子。声音风格大变 由本身的低频偏厚有力 中频不错 高频一般 变成了低频下潜很深但不卖弄 刚刚好 中频、高频趋近绝佳的表现。而且声音也变得更加的干净和明亮 女声更加甜美贴耳。 　　 　　总体来讲： 　　HTC 10低音部分有HTC自己独特的音染 浑厚有力 而最为难得的是在这样的量的低音下中频能有效的分离出来 使得人声表现也很优秀 美中不足的是高音不如前两者那么完美 些许有些吃力（T8ie下表现 Final下就好了很多）。 　　关于杜比耳蜗音效的亮点： 　　 　　1、针对双耳分别去测试 让我想起一句话 来阐述我想说的第一点：世界上没有两片一样的叶子。双手也是一样 双耳更是如此。这样的功能有效的避免了双耳之间因耳道大小不同而出现差异的状况 使得声音完全居中。 　　2、针对不同口味的人群做出了自然的区分 使得调节出来的音效符合自己的口味。 　　3、针对老烧友长时间听音产生的听力衰竭的声音部分有很好的补充。 　　开启调音后声音变得更加立体 声场被强制放大了一些 但声音走向没有变化。 　　相机篇：参数惊艳 算法仍有提升空间 　　相机方面一直是HTC一直想征服 但却一直走得举步维艰的模块。首次搭载UltraPixel相机的HTC One M7亮相以后就引发了一系列的话题 但是400w的像素却令很多用户望而却步。而今HTC 10卷土重来 带来了1200w像素的UltraPixel 让我们来一起看一下详细参数： 　　 　　从参数上我们可以看到光圈提高到f/1.8 这个数值对比M7已经有了较大的提高。 　　 　　从UltraPixel主推的单个像素尺寸方面 HTC 10达到了业界最高的1.55um 完胜其他竞品。 　　 　　 　　加持镭射对焦和光学防抖两大buff单从参数上面确实令人惊艳 我们来看看实际的表现效果 　　室内样张： 　　 　　室外样张： 　　 　　两张样张的表现中规中矩 光线较强的情况下甚至有点拆强人意。 　　暗光与傍晚： 　　 　　 　　而这两张的效果却格外喜人 笔者在拍摄样张的时候也发现了这样的一些细节 比如在拍摄比较细小的枝状物体的时候 相机会默认后方墙面为对焦对象 出现了对不上焦的情况（可利用手动模式解决） 可见拍照算法部分还有很大的提升空间 期待未来升级后的表现。 　　总结： 　　HTC 10更像是总结过往后的一款产品 去掉了吐槽已久的四下巴 电容键回归 将UltraPixel提升至1200w等等改变 虽然配置在当下已经显得有些平庸 但是难能可贵的是HTC这些改变背后表现出的诚意 如果说“若批判不自由则赞美无意义” 那么批判之后应赞美。如果你是一名HTC的老用户正在使用HTC的其他手机 或者是一枚肠粉 我觉得HTC 10是一款好手机 推荐给你购买。但是HTC 10却不是能打得响翻身仗的那款手机 在每况愈下的业绩中不得不让人担忧我们是否可以等到那款翻身旗舰 我们对于HTC寄予了太多的希望和鞭策 愿未来市场除了是能吹者的天下 也能给情怀留一条出路。|http://www.zuinow.com/n1816849.html|2016-05-18
기타|2447741114|sohu_mt|IT|ZHO|2016-05-18 03:56:02|HTC 10：批判不自由 赞美无意义|　　 　　外观篇：宝刀未老 锋芒毕现 　　HTC在工业设计领域一直有着自己对于手机审美的独到见解 在整个手机行业更是独树一帜。HTC 10依然保持高端One系列一贯的金属一体成型的CNC加工工艺 与前代One M9最大的区别就是在于采用了倒角的工艺处理了机身弧形背部与边款衔接 作为工业设计出身的我对于这个设计并没有感到意外 但是这个设计确实使我初见机器概念图的时候就已经迷上这款机器 也在担心万一概念只是概念到最后被砍掉怎么办 但是让人欣喜的是旗舰就是这款产品。 　　 　　这个设计被po出来的时候就有人和我讨论多了这个倒角以后会不会膈手或者割手 但是我拿到真机后得到的体验反馈恰恰是相反的 这样的5mm左右的倒角处理比2mm左右的圆角处理要舒服和自然的多 单手握持时四指第一关节处的压迫感和手掌内侧的压迫感要比M9舒服很多。 　　 　　M9和M10的区别还在于侧边框的设计 虽然从工业美学的角度来看M9的侧边框无论从工艺上还是从设计上都做到了极致 但是这种极致在上市后带来了很多差评 一是整机观感看起来更加厚重（本身就不薄 还搞这一套！）二来侧边手感非常差！（手触摸上去永远是条棱）三来强迫症就是受不了。而10又回归了朴实的处理方式 得益于倒角处理在不影响手感的情况下带来了视觉上更加纤薄的印象（虽然这种设计拍照显得很厚）。 　　 　　另外 细节之处见真功 Sim卡和SD卡卡槽的设置 切实的考虑到了用户应用手机的情景 分别设计在机身边框的两侧 并且放在了靠近顶部的地方 避开了手指可以直接接触的地方 而右侧边框大拇指屈伸范围内分别布置了音量+、音量 – 和坑凹处理过的电源键 让手指可以轻易的就可以接触并区分它们的功能 为这样的设计点赞！ 　　 　　说完了有特色的背部 我们来看一下饱受争议的正脸。 　　说实话 我看到正脸的第一感觉就是为啥指纹识别为什么靠下！不在距离屏幕和边框的边缘 我是强迫症 这样会让我摔手机的 但是使用下来几天以后发现并没有将手机摔掉 而是感觉不到这种问题的存在 个人总结是两个原因带来的 一、我们是竖起来用手机 上下是否对称没有左右是否对称让人敏感；二、这个位置还算舒服 没有带来触感上面的负面反馈。但传感器和前置镜头的位置和设计就不是那么容易让人接受了 如果你恰巧是和我一样的强迫症 恰巧买了白色机器 你恰巧和那几个额头的痣过不去 我劝你还是早点将手机送我吧 因为你早晚会摔掉。（解决方法：1、购买黑色。2、闭眼睛用手机 对于这点如果你想吐槽请参看第一点。） 　　 　　其他一些细节部分： 　　Boomsound扬声器布局做了修改 下方扬声器在边框右下角 而3.5mm耳机插口又被重新移至上方。 　　 　　系统篇：极近原生 不失亮点 　　 　　一开机映入眼帘的就是全新的设置向导界面 这个界面对比之前的老版本的清新了不少但也仅此页面而已 紧接着是几个万年不变的日常设置 增加了指纹识别 其他基本无差别。设置好以后就可以进入系统见到Android6.0和Sense8了 但是给你的第一感觉让我想起了我第一次打开One M7  确实很失望！上一次是陪伴我一个又一个无聊下午的天气动画再也找不到了 这一次恐怕就是Sense再也找不到了 简直让人惋惜。但是上手后感受到的流畅却是前所未有的 或许真的是鱼与熊掌不可兼得吧。 　　 　　极近原生的设置界面： 　　 　　丑陋而实用的相机界面： 　　 　　幸好 标志性的时钟插件还是保留下来了 并且增加了自由主题 这里还是让笔者眼前一亮的。 　　 　　系统界面上对于设置界面和通知栏的布局没有做适当优化确实是令人不满意的地方 但是新的主题模式也使我有了新的乐趣。说完界面我们来讲一下性能 Sense神油是我接触肠粉以来 肠粉们对于HTC手机搭载的系统最好的也是最常用的评价 但是大家对于这个评价往往是从跑分上得来的。笔者一直想说优化和跑分又有什么关系？为了跑分而优化？我觉得是为了使用体验而优化 652版本跑分的正常范围应该在11-13w左右。820版本会在13-15w左右。偶尔跑一下10w 偏低也不能说明什么 放上来只是做一个参考： 　　充电和续航：从未有过的安逸 　　从拿到HTC 10这款机器到成为主力机每天使用感受就两个字“安逸”。这个安逸来自于我重度或者偏重度使用续航仍可以维持一天 只要早晨满电出门一整天都不会担心电量的问题。还有一点就是来自于新的充电技术 当我有急事手机却没有电时 我只要冲几分钟它便可以支撑我打完一个小时电话。下面带来一组安兔兔硬件评测的85%以上电量的评测(评测时忘记了关闭NFC 遗憾)不过仍然得到7279分 我对这个分数处于的阶段并不清楚 而真机在使用的过程当中可以结合各种省电配置 我想这些都是软件给与参考之外的东西。 　　 　　充电方面HTC 10标配一款Quickcharge3.0充电头 这款充电头可以提供更加安全快速的充电体验 实际测试下来亮屏充电从1% 到 42%仅用时30分钟 到实际真正充满也不到2个小时（亮屏） 　　 　　PS: 17:10左右已经充满 此图为后截。 　　音质篇：澎湃音浪 令人难忘 　　在耳机这个圈子也混了很久 结识了很多神人和高手 所以在手机这个圈子很多人都很期待我对手机的音质做一个评测 说实话这让我压力山大 今天就来简单谈谈这门玄学。 　　首先我选择了AK T8ie 、Final VIII、AKG k3003（澳产）来作为本次听音器材。 　　三款耳机在这次测试中也给我们呈现了不一样的声音： 　　AKG K3003： 　　这款耳机应该是大家最熟悉的一款旗舰级入耳耳机了 对于这款耳机也是褒贬不一 但是不可否认的是做工和素质确实一流。 　　 　　在K3003的测试中HTC 10的声音展现出了非常满意的状态 低频饱满有力 中频出色 三频均衡 中正 声音不厚不瘦 展现了非常丰富的声音细节。 　　T8ie： 　　 　　在利用T8ie进行测试的时候 发现HTC 10并不能发挥出T8ie的优秀素质 只能说达到及格的级别 听感如下：T8ie在与10链接后的声音稍厚（t8ie本身就偏厚） 低频和中频表现尚可 人声偏老 高频表现稍微欠佳 有些劈 底噪也稍大。笔者分析造成这样的原因是因为HTC 10尚不能将T8ie完全推开造成的 但是手机能达到这样的状态也是可以接受的。 　　Final Audio heaven VIII 　　 　　这款耳机与10的搭配给我留下了最深刻的印象 给人很意外的感觉就像VIII的靓、柔、甜的裙子给HTC 10这个彪形大汉穿上后 这个大汉居然变成了一个楚楚动人的妹子。声音风格大变 由本身的低频偏厚有力 中频不错 高频一般 变成了低频下潜很深但不卖弄 刚刚好 中频、高频趋近绝佳的表现。而且声音也变得更加的干净和明亮 女声更加甜美贴耳。 　　 　　总体来讲： 　　HTC 10低音部分有HTC自己独特的音染 浑厚有力 而最为难得的是在这样的量的低音下中频能有效的分离出来 使得人声表现也很优秀 美中不足的是高音不如前两者那么完美 些许有些吃力（T8ie下表现 Final下就好了很多）。 　　关于杜比耳蜗音效的亮点： 　　 　　1、针对双耳分别去测试 让我想起一句话 来阐述我想说的第一点：世界上没有两片一样的叶子。双手也是一样 双耳更是如此。这样的功能有效的避免了双耳之间因耳道大小不同而出现差异的状况 使得声音完全居中。 　　2、针对不同口味的人群做出了自然的区分 使得调节出来的音效符合自己的口味。 　　3、针对老烧友长时间听音产生的听力衰竭的声音部分有很好的补充。 　　开启调音后声音变得更加立体 声场被强制放大了一些 但声音走向没有变化。 　　相机篇：参数惊艳 算法仍有提升空间 　　相机方面一直是HTC一直想征服 但却一直走得举步维艰的模块。首次搭载UltraPixel相机的HTC One M7亮相以后就引发了一系列的话题 但是400w的像素却令很多用户望而却步。而今HTC 10卷土重来 带来了1200w像素的UltraPixel 让我们来一起看一下详细参数： 　　 　　从参数上我们可以看到光圈提高到f/1.8 这个数值对比M7已经有了较大的提高。 　　 　　从UltraPixel主推的单个像素尺寸方面 HTC 10达到了业界最高的1.55um 完胜其他竞品。 　　 　　 　　加持镭射对焦和光学防抖两大buff单从参数上面确实令人惊艳 我们来看看实际的表现效果 　　室内样张： 　　 　　室外样张： 　　 　　两张样张的表现中规中矩 光线较强的情况下甚至有点拆强人意。 　　暗光与傍晚： 　　 　　 　　而这两张的效果却格外喜人 笔者在拍摄样张的时候也发现了这样的一些细节 比如在拍摄比较细小的枝状物体的时候 相机会默认后方墙面为对焦对象 出现了对不上焦的情况（可利用手动模式解决） 可见拍照算法部分还有很大的提升空间 期待未来升级后的表现。 　　总结： 　　HTC 10更像是总结过往后的一款产品 去掉了吐槽已久的四下巴 电容键回归 将UltraPixel提升至1200w等等改变 虽然配置在当下已经显得有些平庸 但是难能可贵的是HTC这些改变背后表现出的诚意 如果说“若批判不自由则赞美无意义” 那么批判之后应赞美。如果你是一名HTC的老用户正在使用HTC的其他手机 或者是一枚肠粉 我觉得HTC 10是一款好手机 推荐给你购买。但是HTC 10却不是能打得响翻身仗的那款手机 在每况愈下的业绩中不得不让人担忧我们是否可以等到那款翻身旗舰 我们对于HTC寄予了太多的希望和鞭策 愿未来市场除了是能吹者的天下 也能给情怀留一条出路。|http://mt.sohu.com/20160518/n450025801.shtml|2016-05-18
기타|2447765893|haixiaol|IT科技 最新更新|ZHO|2016-05-18 04:33:01|HTC 10：批判不自由 贊美無意義|　　 　　外觀篇：寶刀未老 鋒芒畢現 　　HTC在工業設計領域一直有著自己對于手機審美的獨到見解 在整個手機行業更是獨樹一幟。HTC 10依然保持高端One系列一貫的金屬一體成型的CNC加工工藝 與前代One M9最大的區別就是在于采用了倒角的工藝處理了機身弧形背部與邊款銜接 作為工業設計出身的我對于這個設計并沒有感到意外 但是這個設計確實使我初見機器概念圖的時候就已經迷上這款機器 也在擔心萬一概念只是概念到最后被砍掉怎么辦 但是讓人欣喜的是旗艦就是這款產品。 　　 　　這個設計被po出來的時候就有人和我討論多了這個倒角以后會不會膈手或者割手 但是我拿到真機后得到的體驗反饋恰恰是相反的 這樣的5mm左右的倒角處理比2mm左右的圓角處理要舒服和自然的多 單手握持時四指第一關節處的壓迫感和手掌內側的壓迫感要比M9舒服很多。 　　 　　M9和M10的區別還在于側邊框的設計 雖然從工業美學的角度來看M9的側邊框無論從工藝上還是從設計上都做到了極致 但是這種極致在上市后帶來了很多差評 一是整機觀感看起來更加厚重（本身就不薄 還搞這一套！）二來側邊手感非常差！（手觸摸上去永遠是條棱）三來強迫癥就是受不了。而10又回歸了樸實的處理方式 得益于倒角處理在不影響手感的情況下帶來了視覺上更加纖薄的印象（雖然這種設計拍照顯得很厚）。 　　 　　另外 細節之處見真功 Sim卡和SD卡卡槽的設置 切實的考慮到了用戶應用手機的情景 分別設計在機身邊框的兩側 并且放在了靠近頂部的地方 避開了手指可以直接接觸的地方 而右側邊框大拇指屈伸范圍內分別布置了音量+、音量 – 和坑凹處理過的電源鍵 讓手指可以輕易的就可以接觸并區分它們的功能 為這樣的設計點贊！ 　　 　　說完了有特色的背部 我們來看一下飽受爭議的正臉。 　　說實話 我看到正臉的第一感覺就是為啥指紋識別為什么靠下！不在距離熒幕和邊框的邊緣 我是強迫癥 這樣會讓我摔手機的 但是使用下來幾天以后發現并沒有將手機摔掉 而是感覺不到這種問題的存在 個人總結是兩個原因帶來的 一、我們是豎起來用手機 上下是否對稱沒有左右是否對稱讓人敏感；二、這個位置還算舒服 沒有帶來觸感上面的負面反饋。但傳感器和前置鏡頭的位置和設計就不是那么容易讓人接受了 如果你恰巧是和我一樣的強迫癥 恰巧買了白色機器 你恰巧和那幾個額頭的痣過不去 我勸你還是早點將手機送我吧 因為你早晚會摔掉。（解決方法：1、購買黑色。2、閉眼睛用手機 對于這點如果你想吐槽請參看第一點。） 　　 　　其他一些細節部分： 　　Boomsound揚聲器布局做了修改 下方揚聲器在邊框右下角 而3.5mm耳機插口又被重新移至上方。 　　 　　系統篇：極近原生 不失亮點 　　 　　一開機映入眼簾的就是全新的設置向導界面 這個界面對比之前的老版本的清新了不少但也僅此頁面而已 緊接著是幾個萬年不變的日常設置 增加了指紋識別 其他基本無差別。設置好以后就可以進入系統見到Android6.0和Sense8了 但是給你的第一感覺讓我想起了我第一次打開One M7  確實很失望！上一次是陪伴我一個又一個無聊下午的天氣動畫再也找不到了 這一次恐怕就是Sense再也找不到了 簡直讓人惋惜。但是上手后感受到的流暢卻是前所未有的 或許真的是魚與熊掌不可兼得吧。 　　 　　極近原生的設置界面： 　　 　　丑陋而實用的相機界面： 　　 　　幸好 標志性的時鐘插件還是保留下來了 并且增加了自由主題 這里還是讓筆者眼前一亮的。 　　 　　系統界面上對于設置界面和訊息欄的布局沒有做適當優化確實是令人不滿意的地方 但是新的主題模式也使我有了新的樂趣。說完界面我們來講一下性能 Sense神油是我接觸腸粉以來 腸粉們對于HTC手機搭載的系統最好的也是最常用的評價 但是大家對于這個評價往往是從跑分上得來的。筆者一直想說優化和跑分又有什么關系？為了跑分而優化？我覺得是為了使用體驗而優化 652版本跑分的正常范圍應該在11-13w左右。820版本會在13-15w左右。偶爾跑一下10w 偏低也不能說明什么 放上來只是做一個參考： 　　充電和續航：從未有過的安逸 　　從拿到HTC 10這款機器到成為主力機每天使用感受就兩個字“安逸”。這個安逸來自于我重度或者偏重度使用續航仍可以維持一天 只要早晨滿電出門一整天都不會擔心電量的問題。還有一點就是來自于新的充電技術 當我有急事手機卻沒有電時 我只要沖幾分鐘它便可以支撐我打完一個小時電話。下面帶來一組安兔兔硬件評測的85%以上電量的評測(評測時忘記了關閉NFC 遺憾)不過仍然得到7279分 我對這個分數處于的階段并不清楚 而真機在使用的過程當中可以結合各種省電配置 我想這些都是軟體給與參考之外的東西。 　　 　　充電方面HTC 10標配一款Quickcharge3.0充電頭 這款充電頭可以提供更加安全快速的充電體驗 實際測試下來亮屏充電從1% 到 42%僅用時30分鐘 到實際真正充滿也不到2個小時（亮屏） 　　 　　PS: 17:10左右已經充滿 此圖為后截。 　　音質篇：澎湃音浪 令人難忘 　　在耳機這個圈子也混了很久 結識了很多神人和高手 所以在手機這個圈子很多人都很期待我對手機的音質做一個評測 說實話這讓我壓力山大 今天就來簡單談談這門玄學。 　　首先我選擇了AK T8ie 、Final VIII、AKG k3003（澳產）來作為本次聽音器材。 　　三款耳機在這次測試中也給我們呈現了不一樣的聲音： 　　AKG K3003： 　　這款耳機應該是大家最熟悉的一款旗艦級入耳耳機了 對于這款耳機也是褒貶不一 但是不可否認的是做工和貭素確實一流。 　　 　　在K3003的測試中HTC 10的聲音展現出了非常滿意的狀態 低頻飽滿有力 中頻出色 三頻均衡 中正 聲音不厚不瘦 展現了非常豐富的聲音細節。 　　T8ie： 　　 　　在利用T8ie進行測試的時候 發現HTC 10并不能發揮出T8ie的優秀貭素 只能說達到及格的級別 聽感如下：T8ie在與10鏈接后的聲音稍厚（t8ie本身就偏厚） 低頻和中頻表現尚可 人聲偏老 高頻表現稍微欠佳 有些劈 底噪也稍大。筆者分析造成這樣的原因是因為HTC 10尚不能將T8ie完全推開造成的 但是手機能達到這樣的狀態也是可以接受的。 　　Final Audio heaven VIII 　　 　　這款耳機與10的搭配給我留下了最深刻的印象 給人很意外的感覺就像VIII的靚、柔、甜的裙子給HTC 10這個彪形大漢穿上后 這個大漢居然變成了一個楚楚動人的妹子。聲音風格大變 由本身的低頻偏厚有力 中頻不錯 高頻一般 變成了低頻下潛很深但不賣弄 剛剛好 中頻、高頻趨近絕佳的表現。而且聲音也變得更加的干凈和明亮 女聲更加甜美貼耳。 　　 　　總體來講： 　　HTC 10低音部分有HTC自己獨特的音染 渾厚有力 而最為難得的是在這樣的量的低音下中頻能有效的分離出來 使得人聲表現也很優秀 美中不足的是高音不如前兩者那么完美 些許有些吃力（T8ie下表現 Final下就好了很多）。 　　關于杜比耳蝸音效的亮點： 　　 　　1、針對雙耳分別去測試 讓我想起一句話 來闡述我想說的第一點：世界上沒有兩片一樣的葉子。雙手也是一樣 雙耳更是如此。這樣的功能有效的避免了雙耳之間因耳道大小不同而出現差異的狀況 使得聲音完全居中。 　　2、針對不同口味的人群做出了自然的區分 使得調節出來的音效符合自己的口味。 　　3、針對老燒友長時間聽音產生的聽力衰竭的聲音部分有很好的補充。 　　開啟調音后聲音變得更加立體 聲場被強制放大了一些 但聲音走向沒有變化。 　　相機篇：參數驚艷 算法仍有提升空間 　　相機方面一直是HTC一直想征服 但卻一直走得舉步維艱的模塊。首次搭載UltraPixel相機的HTC One M7亮相以后就引發了一系列的話題 但是400w的像素卻令很多用戶望而卻步。而今HTC 10卷土重來 帶來了1200w像素的UltraPixel 讓我們來一起看一下詳細參數： 　　 　　從參數上我們可以看到光圈提高到f/1.8 這個數值對比M7已經有了較大的提高。 　　 　　從UltraPixel主推的單個像素尺寸方面 HTC 10達到了業界最高的1.55um 完勝其他競品。 　　 　　 　　加持鐳射對焦和光學防抖兩大buff單從參數上面確實令人驚艷 我們來看看實際的表現效果 　　室內樣張： 　　 　　室外樣張： 　　 　　兩張樣張的表現中規中矩 光線較強的情況下甚至有點拆強人意。 　　暗光與傍晚： 　　 　　 　　而這兩張的效果卻格外喜人 筆者在拍攝樣張的時候也發現了這樣的一些細節 比如在拍攝比較細小的枝狀物體的時候 相機會默認后方墻面為對焦對象 出現了對不上焦的情況（可利用手動模式解決） 可見拍照算法部分還有很大的提升空間 期待未來升級后的表現。 　　總結： 　　HTC 10更像是總結過往后的一款產品 去掉了吐槽已久的四下巴 電容鍵回歸 將UltraPixel提升至1200w等等改變 雖然配置在當下已經顯得有些平庸 但是難能可貴的是HTC這些改變背后表現出的誠意 如果說“若批判不自由則贊美無意義” 那么批判之后應贊美。如果你是一名HTC的老用戶正在使用HTC的其他手機 或者是一枚腸粉 我覺得HTC 10是一款好手機 推薦給你購買。但是HTC 10卻不是能打得響翻身仗的那款手機 在每況愈下的業績中不得不讓人擔憂我們是否可以等到那款翻身旗艦 我們對于HTC寄予了太多的希望和鞭策 愿未來市場除了是能吹者的天下 也能給情懷留一條出路。|http://www.haixiaol.com/n1814312.html|2016-05-18
기타|2447780022|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-18 04:55:02|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=53&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-18
기타|2447816702|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-18 05:53:01|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=54&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-18
기타|2448027239|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-18 09:38:02|2016年04月14日 发表了口碑|来自：手机汽车之家  2016年04月14日 发表了口碑  口碑    《不是一般的省油 跟1.6排量的一个油耗 保养便宜 省心省力！》           【最满意的一点】省油 不是一般的省油 100块大洋 跑200 公里很容易 保养也便宜 在4s小保一次300多块 换的是麦戈龙的半合成！用着还可以！【最不满意的一点】车漆太薄了 减震略硬 主副驾驶都有异响 比较烦人 就是找不到原因！高速给人信心略有不足！其他还好！【空间】空间相当的大 后排3个胖子毫无压力！后备箱我总装货 装的满满的 【动力】起步比较肉 不过过了60以后还可以 够用而已 高速超车还是比较有信心。挂上s档 在高速 感觉点油门嗖嗖的 或许3000转以后才会有动力！【操控】转向精准 方向盘比较小 操控如鱼得水！就是车头的位置总看不好！【油耗】相当省油.跟家里另台1.6的k3一个油后 甚至更省油！高速神器！【舒适性】座椅宽大 挺舒服 但是时间久了腰比较累 可能没有支撑的作用！【外观】外观大气 前脸很唬人 比较霸气！【内饰】内饰做工精致 仪表台软性材质 科技感比较好！【性价比】物有所值！性价比还是比较高的。【为什么最终选择这款车？】当初看了凯美瑞 价格优惠比较大 也比较皮实 但是因为要改款 而且4速是最不能接受的！韩系 美系不再考虑范围之内 大众哥俩因为价格略贵 也pass了 不过个人还是挺喜欢这哥俩的 最后因为9代雅阁刚换代不久 而且价格也比较吸引人 再加上本田的车皮实耐用 省心 省油 后期的保养也便宜 就选择了丐版的雅9！【其他描述】雅9快2年了 没出现过什么问题 比较省心 不后悔拥有！|http://k.autohome.com.cn/spec/18279/view_1070627_1.html?st=197&piap=0 78 0 0 2 0 0 0 0 0 1#20160414|2016-05-18
기타|2448027675|Autohome_review|혼다 어코드(雅阁)|ZHO|2016-05-18 09:38:03|2016年05月09日 发表了口碑|来自：手机汽车之家  2016年05月09日 发表了口碑  口碑    《你是我最重要的决定！附上全车亚光黑效果图！》             【最满意的一点】一、大 真大 小雅的身体里不是一般的大 开习惯小雅在开盆友的卡罗拉感觉腿都伸不开 本人1.83～～～二、动力 都说2.0的动力拉小雅的身体有点吃力 可我感觉很好 主要是舍不舍得踩 等红灯基本上都是我第一个出去 （喷子们别说什么别的车懒得踩油门哈）总得来说动力对我足够用了。三、油耗 小雅的油耗不高 小弟我住在县级市 离市里30公里 一个月也进不几趟城 其余的道路状况基本没有堵车畅通的很9个油【最不满意的一点】不难意的地方嘛 中控的异响 不过本人没音乐不开车 所以忽略。A柱的视线不好这点很重要。还有就是用u盘听歌有时候会显示未连接 只需要把u盘拔了重新插上就好了。【空间】大 真大 真心的大 在车里自由的折腾了 你们懂得！【动力】 只要舍得踩油门动力绝对可以满足你想要的一切！【操控】 没开过什么好车 雅阁的方向感很好 悬架支撑的还算可以。【油耗】基本上保持在8 9个  本人脚重。【舒适性】提速轻盈 走坏路也感觉不出太颠 一直也没坐在后面过但是坐在后面的都说真舒服 钱不白花！【外观】小雅的霸气是无人能敌的（在我心里）大龅牙日行灯真是越看越喜欢。【内饰】内饰感觉很简洁 没有改装大屏喜欢原汁原味 用料上也很厚道 就是小异响有点瑕疵。【性价比】配置很好 最低配想要的也都齐全 价格的话没在意那么多因为是分期还多少也没太在意。【为什么最终选择这款车？】选车真是痛苦的事情 当时是看了紧凑型的车 卡罗拉 雷凌  捷达 桑塔纳 朗逸 朗行 k3 朗动 轩逸 哈佛H6 长安CS75 这些都是我能接受了的车型  经过一一筛选最后只剩下了雷凌跟轩逸 （详情请看提车作业） 至于最后为什么买了小雅完全是预料之外的情况 一年的时间让我对小雅是越来越喜欢 半一年的时间也让我对它进行了改变～【其他描述】|http://k.autohome.com.cn/spec/22135/view_1106334_1.html?st=45&piap=0 78 0 0 2 0 0 0 0 0 1#20160509|2016-05-18
기타|2448401406|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-18 13:22:33|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=55&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-18
各大媒体|2448423697|gmw|滚动读报|ZHO|2016-05-18 13:36:01|改变自己 由内到外 新k3散发全新风采|"url:http://epaper.tianjinwe.com/tjrb/tjrb/2016-05/18/content_*******.htm|id:0健身风潮近两年热度不减 人们开始通过运动来塑造自己的全新形象。说到新形象 小编要推荐一款由内到外都进行了全面升级 带来全新风采的车型——东风悦达起亚新k3。全新升级的新k3采用年轻、干练、高端大气的前后脸设计 使整体造型更为稳重、大气。改变 最终要落到内芯。新k3拥有1.4t及1.6l两种动力总成 兼具高性能、高输出与耐久性的优势。现在购买新k3可享受24期“0利息0手续费”信贷政策（24期贷款0利息0手续费仅限银行政策） 以及“0购置税”的惊喜购车优惠。你做好准备 和新k3一起去改变自己了吗？"|http://news.gmw.cn/newspaper/2016-05/18/content_112541948.htm|2016-05-18
기타|2448509930|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-18 14:28:52|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=57&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-18
기타|2448538461|Autohome_review|잉랑GT(英朗)|ZHO|2016-05-18 14:45:03|2016年05月14日 发表了口碑|"2016年05月14日 发表了口碑  口碑    《全新英朗买的值！推荐》           本人今年本命年 24了还没有个对象 以前上学的时候觉得工作了以后找对象 工作了发现根本不是那一回事 工作了2年多 也没攒下多少钱 又到了结婚的年纪 人丑读书还不多 家里有点着急了 给我买了一辆车 让我这样看起来好找对象。（聊得有点多了 见谅！） 我是15年的45月份就开始关注汽车 当时看的也比较多 一开始在考虑国产车 后来让朋友同学同事说的 买国产没大谱 又开始考虑合资车 10w多的车 就比较多了 科鲁兹 福克斯 福睿斯 朗动 名图 k3 世嘉 卡罗拉 雷凌 宝来 朗逸 天天看咱们汽车之家的图片和朋友们的评价 这些车也没有什么可多说的了 就像看女人一样 能入你眼的 你才会去研究了解 当时我就筛去了一些 留下科鲁兹 福克斯 福睿斯 和朗逸了 当然还有全新英朗 先从外形来说 全新英朗我觉得最漂亮 再就是科鲁兹了 福克斯 朗逸 卡罗拉。当时就想着就从这几款车里选吧 有空的时候去4s店试驾一下 什么的。科鲁兹这款车 挺好的 新科操控没得说 很棒 就是车头太小了 感觉和新赛欧的似的 经典款的 还不错 但是我比较纠结两个地方 一个内饰的按键太多 显得很乱 再一个就是他的发动机动静 感觉和拖拉机似的 我把科鲁兹就给筛去了 福克斯 朗逸 卡罗拉 感觉都不错的 优缺点不说了 但我说个全新英朗最实用的优点就是 后排空间要比这几款车都大 还有吸人眼球的LED日行灯 实用加时尚 最后就在15年的10月2号 在车展上定了车 11月低 才提的车。【最满意的一点】油耗是我没真想到的 空间 外形。【最不满意的一点】最不满意的就是夜间的时候 车内门碗没有小灯 夜间下车找不到把手。还有就是开车门 就亮内饰灯 不管是白天黑夜。【空间】后排很舒适 朋友喜欢后排（同级别车）【动力】动力也不错 我6.5个油 当然也不是慢腾腾的 我也喜欢刺激 上下班太堵 所以经常超车 舍得给油 动力也是可以的。【操控】还不错吧 没有长时间驾驶过其他车 舒适型的吧【油耗】现在6000公里 我现在才发贴 因为我自己都有点不相信 但是我要告诉大家【舒适性】很好 独立悬挂很舒适【外观】亮点就是LED日行灯了【内饰】还算可以 还没换中控屏 暂时用的收音机【性价比】很高了【其它描述】刚刚提车的时候 不知道是不是自己的驾驶问题 还是路面问题 老是感觉 车快满载在过坑的时候车屁股左右晃动 而且乘坐的人都能感觉到 有懂朋友吗?能给解释一下不？【为什么最终选择这款车】第一外形 第二空间 第三优惠了1.7w说了很多 不知道现在还有没有人关注全新英朗 新车这么多 现在也出2016款的了 更值得选购了 油耗真的只有自己开了 才会相信 证明车的油耗 我可以以后追加的 考虑这款车的朋友可以留言给我。谢谢大家支持！（手机拍的照片太大|没法发图认证车主了 见谅 拍的图片很多就一个能上传）"|http://k.autohome.com.cn/spec/21677/view_1113219_1.html?st=58&piap=0 982 0 0 2 0 0 0 0 0 1#20160514|2016-05-18
기타|2448687305|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-18 16:09:02|2016年05月09日 发表了口碑|"来自：手机汽车之家  2016年05月09日 发表了口碑  口碑   《动力强劲 省油 提速快 噪音小》           【最满意的一点】低油耗 动力足 【最不满意的一点】车身接缝太大。【空间】家用刚好【动力】提速超车很快 【操控】转向非常精确和灵敏 【油耗】油耗超乎我的想象【舒适性】整体舒适还不错 要有后独立悬架就好了【外观】外观是我最喜欢的 犀利前卫时尚【内饰】内饰这个价钱的车可以了【性价比】就是这个价位没有esp【为什么最终选择这款车？】看了别克新英朗 现代朗动 起亚k3.日产轩逸 朗逸  别克英朗的日行灯是大爱可是尾部太小气了 整个就是加大版的凯越记录仪朗动动力和外观各方面都挺满意 就是车身和头部太短了直接pass 日产轩逸差点就定 就是缩小版的小天籁 挺喜欢 后来听朋友说烧机油。也无奈pass|然后就是k3前脸和尾部都满意 就是日行灯太单调不喜欢最后就是朗逸 简直就是神车 后来出来了尾气门事件 pass||最后看到卡罗拉各种喜【其他描述】整体还不错 建议购买"|http://k.autohome.com.cn/spec/18889/view_1105663_1.html?st=69&piap=0 526 0 0 2 0 0 0 0 0 1#20160509|2016-05-18
기타|2448687420|Autohome_review|뉴 코롤라(卡罗拉)|ZHO|2016-05-18 16:09:02|2016年05月13日 发表了口碑|来自：手机汽车之家  2016年05月13日 发表了口碑  口碑   《油耗低 空间大 动力足 外表炫酷 喜欢的没话说》   【最满意的一点】最喜欢的就是空间和动力方面了 空间没的说大家都公认的大有人说动力只是一般我试过一车五人八百多斤  因为像我姑啥的比较胖当时我都心疼车新车啊  但是起步路上跑啥的动力绰绰有余 也可能是我新手的原因吧没来过啥好车这动力已经非常满足了 只能说没有动力差的车只要舍得踩油 卡卡的动力还是很好的【最不满意的一点】离合有点高  刚开始不是很适应  后来慢慢的摸索习惯了开着很顺手  因为资金方面买的手动低配没有发动机安全锁比较遗憾 跟中配对比了一下仪表盘视觉方面还是差了点 另外不带座椅升降感觉档次低了不少 但是一分钱一分货嘛 总体感觉还是很不错的 值得一说的是后视镜调到正常驾驶的角度看不到底部 家是农村的平时避免不了走窄路偶尔倒车看不到地面哪里有沟还得来回调角度感觉挺不方便的 以前练车时候根本没注意到这个问题【空间】卡卡的内部空间那真是没的说尤其后排空间三个稍微偏胖的成年人不觉得拥挤这一点家里人比较满意毕竟除了我比较瘦以外家里人都是有点偏胖型的都是170斤往上的那种他们都不嫌弃挤我当然更是没话说喽【动力】动力方面还是很不错的刚提车那会开车非常小心毕竟还在实习期嘛一直都是用怠速起步也不觉得慢后来慢慢的摸索清楚了就有点不太满足了起步开始踩油门不得不说只要舍得给油动力很不错路上正常行驶三档超车动力绰绰有余非常给力【操控】指向非常精准属于指哪打哪那种很满意路面反馈很好 农村的路面坑坑洼洼的很难走 但是卡卡悬挂设计的不错颠簸很化解的很轻微不会产生颠簸的难受那种感觉 每次走在这种路面我都把颠簸当成按摩了 哈哈【油耗】预期新手能跑出8.0左右油耗就不错了没想到能跑出7.1油耗  满意的没话说【舒适性】座椅舒适度还是不错的我比较瘦坐在驾驶座上空间余量比较大估计是按照成年人的体型设计的吧 不过噪音方面感觉还是有提神空间的尤其小石子打在底盘上声音确实有点烦人虽然开车喜欢放音乐但是毕竟不是所有人都喜欢边开车边听歌的吧【外观】外观是我最喜欢的地方尤其是前脸车灯喜欢的无药可救了选择卡卡很大一部分原因就是外观了如果说我有病那卡卡就是药【内饰】中控台用的软材料底部才是硬塑料设计的不错【性价比】配置方面感觉发动机防盗应该标配  安全嘛【为什么最终选择这款车？】从家里人说买车到订车看了一个月的汽车之家刚开始打算十万以内落地关注了景逸x5 比亚迪s6后来想想国产车实在有点让人心寒转战合资车朗动  k3韩国车配置要高点便宜点但是实在没看好设计方面 可能当时也是倾心卡罗拉的原因吧  想来想去一咬牙就选卡卡了  丑了个时间试驾都省了直接订车 车是从老爷子的一个朋友那里定的 所以没法讲价说了个最低价就交钱了  等了大约得半个月  就提车了【其他描述】|http://k.autohome.com.cn/spec/18889/view_1112492_1.html?st=23&piap=0 526 0 0 2 0 0 0 0 0 1#20160513|2016-05-18
